
module MULT(A, B, P);

    //ports
    input [71:0] A;
    input [40:0] B;

    output [112:0] P;


    //wire names
    wire stage0_r0_c0;
    wire stage0_r0_c1;
    wire stage0_r1_c0;
    wire stage0_r0_c2;
    wire stage0_r1_c1;
    wire stage0_r2_c0;
    wire stage0_r0_c3;
    wire stage0_r1_c2;
    wire stage0_r2_c1;
    wire stage0_r3_c0;
    wire stage0_r0_c4;
    wire stage0_r1_c3;
    wire stage0_r2_c2;
    wire stage0_r3_c1;
    wire stage0_r4_c0;
    wire stage0_r0_c5;
    wire stage0_r1_c4;
    wire stage0_r2_c3;
    wire stage0_r3_c2;
    wire stage0_r4_c1;
    wire stage0_r5_c0;
    wire stage0_r0_c6;
    wire stage0_r1_c5;
    wire stage0_r2_c4;
    wire stage0_r3_c3;
    wire stage0_r4_c2;
    wire stage0_r5_c1;
    wire stage0_r6_c0;
    wire stage0_r0_c7;
    wire stage0_r1_c6;
    wire stage0_r2_c5;
    wire stage0_r3_c4;
    wire stage0_r4_c3;
    wire stage0_r5_c2;
    wire stage0_r6_c1;
    wire stage0_r7_c0;
    wire stage0_r0_c8;
    wire stage0_r1_c7;
    wire stage0_r2_c6;
    wire stage0_r3_c5;
    wire stage0_r4_c4;
    wire stage0_r5_c3;
    wire stage0_r6_c2;
    wire stage0_r7_c1;
    wire stage0_r8_c0;
    wire stage0_r0_c9;
    wire stage0_r1_c8;
    wire stage0_r2_c7;
    wire stage0_r3_c6;
    wire stage0_r4_c5;
    wire stage0_r5_c4;
    wire stage0_r6_c3;
    wire stage0_r7_c2;
    wire stage0_r8_c1;
    wire stage0_r9_c0;
    wire stage0_r0_c10;
    wire stage0_r1_c9;
    wire stage0_r2_c8;
    wire stage0_r3_c7;
    wire stage0_r4_c6;
    wire stage0_r5_c5;
    wire stage0_r6_c4;
    wire stage0_r7_c3;
    wire stage0_r8_c2;
    wire stage0_r9_c1;
    wire stage0_r10_c0;
    wire stage0_r0_c11;
    wire stage0_r1_c10;
    wire stage0_r2_c9;
    wire stage0_r3_c8;
    wire stage0_r4_c7;
    wire stage0_r5_c6;
    wire stage0_r6_c5;
    wire stage0_r7_c4;
    wire stage0_r8_c3;
    wire stage0_r9_c2;
    wire stage0_r10_c1;
    wire stage0_r11_c0;
    wire stage0_r0_c12;
    wire stage0_r1_c11;
    wire stage0_r2_c10;
    wire stage0_r3_c9;
    wire stage0_r4_c8;
    wire stage0_r5_c7;
    wire stage0_r6_c6;
    wire stage0_r7_c5;
    wire stage0_r8_c4;
    wire stage0_r9_c3;
    wire stage0_r10_c2;
    wire stage0_r11_c1;
    wire stage0_r12_c0;
    wire stage0_r0_c13;
    wire stage0_r1_c12;
    wire stage0_r2_c11;
    wire stage0_r3_c10;
    wire stage0_r4_c9;
    wire stage0_r5_c8;
    wire stage0_r6_c7;
    wire stage0_r7_c6;
    wire stage0_r8_c5;
    wire stage0_r9_c4;
    wire stage0_r10_c3;
    wire stage0_r11_c2;
    wire stage0_r12_c1;
    wire stage0_r13_c0;
    wire stage0_r0_c14;
    wire stage0_r1_c13;
    wire stage0_r2_c12;
    wire stage0_r3_c11;
    wire stage0_r4_c10;
    wire stage0_r5_c9;
    wire stage0_r6_c8;
    wire stage0_r7_c7;
    wire stage0_r8_c6;
    wire stage0_r9_c5;
    wire stage0_r10_c4;
    wire stage0_r11_c3;
    wire stage0_r12_c2;
    wire stage0_r13_c1;
    wire stage0_r14_c0;
    wire stage0_r0_c15;
    wire stage0_r1_c14;
    wire stage0_r2_c13;
    wire stage0_r3_c12;
    wire stage0_r4_c11;
    wire stage0_r5_c10;
    wire stage0_r6_c9;
    wire stage0_r7_c8;
    wire stage0_r8_c7;
    wire stage0_r9_c6;
    wire stage0_r10_c5;
    wire stage0_r11_c4;
    wire stage0_r12_c3;
    wire stage0_r13_c2;
    wire stage0_r14_c1;
    wire stage0_r15_c0;
    wire stage0_r0_c16;
    wire stage0_r1_c15;
    wire stage0_r2_c14;
    wire stage0_r3_c13;
    wire stage0_r4_c12;
    wire stage0_r5_c11;
    wire stage0_r6_c10;
    wire stage0_r7_c9;
    wire stage0_r8_c8;
    wire stage0_r9_c7;
    wire stage0_r10_c6;
    wire stage0_r11_c5;
    wire stage0_r12_c4;
    wire stage0_r13_c3;
    wire stage0_r14_c2;
    wire stage0_r15_c1;
    wire stage0_r16_c0;
    wire stage0_r0_c17;
    wire stage0_r1_c16;
    wire stage0_r2_c15;
    wire stage0_r3_c14;
    wire stage0_r4_c13;
    wire stage0_r5_c12;
    wire stage0_r6_c11;
    wire stage0_r7_c10;
    wire stage0_r8_c9;
    wire stage0_r9_c8;
    wire stage0_r10_c7;
    wire stage0_r11_c6;
    wire stage0_r12_c5;
    wire stage0_r13_c4;
    wire stage0_r14_c3;
    wire stage0_r15_c2;
    wire stage0_r16_c1;
    wire stage0_r17_c0;
    wire stage0_r0_c18;
    wire stage0_r1_c17;
    wire stage0_r2_c16;
    wire stage0_r3_c15;
    wire stage0_r4_c14;
    wire stage0_r5_c13;
    wire stage0_r6_c12;
    wire stage0_r7_c11;
    wire stage0_r8_c10;
    wire stage0_r9_c9;
    wire stage0_r10_c8;
    wire stage0_r11_c7;
    wire stage0_r12_c6;
    wire stage0_r13_c5;
    wire stage0_r14_c4;
    wire stage0_r15_c3;
    wire stage0_r16_c2;
    wire stage0_r17_c1;
    wire stage0_r18_c0;
    wire stage0_r0_c19;
    wire stage0_r1_c18;
    wire stage0_r2_c17;
    wire stage0_r3_c16;
    wire stage0_r4_c15;
    wire stage0_r5_c14;
    wire stage0_r6_c13;
    wire stage0_r7_c12;
    wire stage0_r8_c11;
    wire stage0_r9_c10;
    wire stage0_r10_c9;
    wire stage0_r11_c8;
    wire stage0_r12_c7;
    wire stage0_r13_c6;
    wire stage0_r14_c5;
    wire stage0_r15_c4;
    wire stage0_r16_c3;
    wire stage0_r17_c2;
    wire stage0_r18_c1;
    wire stage0_r19_c0;
    wire stage0_r0_c20;
    wire stage0_r1_c19;
    wire stage0_r2_c18;
    wire stage0_r3_c17;
    wire stage0_r4_c16;
    wire stage0_r5_c15;
    wire stage0_r6_c14;
    wire stage0_r7_c13;
    wire stage0_r8_c12;
    wire stage0_r9_c11;
    wire stage0_r10_c10;
    wire stage0_r11_c9;
    wire stage0_r12_c8;
    wire stage0_r13_c7;
    wire stage0_r14_c6;
    wire stage0_r15_c5;
    wire stage0_r16_c4;
    wire stage0_r17_c3;
    wire stage0_r18_c2;
    wire stage0_r19_c1;
    wire stage0_r20_c0;
    wire stage0_r0_c21;
    wire stage0_r1_c20;
    wire stage0_r2_c19;
    wire stage0_r3_c18;
    wire stage0_r4_c17;
    wire stage0_r5_c16;
    wire stage0_r6_c15;
    wire stage0_r7_c14;
    wire stage0_r8_c13;
    wire stage0_r9_c12;
    wire stage0_r10_c11;
    wire stage0_r11_c10;
    wire stage0_r12_c9;
    wire stage0_r13_c8;
    wire stage0_r14_c7;
    wire stage0_r15_c6;
    wire stage0_r16_c5;
    wire stage0_r17_c4;
    wire stage0_r18_c3;
    wire stage0_r19_c2;
    wire stage0_r20_c1;
    wire stage0_r21_c0;
    wire stage0_r0_c22;
    wire stage0_r1_c21;
    wire stage0_r2_c20;
    wire stage0_r3_c19;
    wire stage0_r4_c18;
    wire stage0_r5_c17;
    wire stage0_r6_c16;
    wire stage0_r7_c15;
    wire stage0_r8_c14;
    wire stage0_r9_c13;
    wire stage0_r10_c12;
    wire stage0_r11_c11;
    wire stage0_r12_c10;
    wire stage0_r13_c9;
    wire stage0_r14_c8;
    wire stage0_r15_c7;
    wire stage0_r16_c6;
    wire stage0_r17_c5;
    wire stage0_r18_c4;
    wire stage0_r19_c3;
    wire stage0_r20_c2;
    wire stage0_r21_c1;
    wire stage0_r22_c0;
    wire stage0_r0_c23;
    wire stage0_r1_c22;
    wire stage0_r2_c21;
    wire stage0_r3_c20;
    wire stage0_r4_c19;
    wire stage0_r5_c18;
    wire stage0_r6_c17;
    wire stage0_r7_c16;
    wire stage0_r8_c15;
    wire stage0_r9_c14;
    wire stage0_r10_c13;
    wire stage0_r11_c12;
    wire stage0_r12_c11;
    wire stage0_r13_c10;
    wire stage0_r14_c9;
    wire stage0_r15_c8;
    wire stage0_r16_c7;
    wire stage0_r17_c6;
    wire stage0_r18_c5;
    wire stage0_r19_c4;
    wire stage0_r20_c3;
    wire stage0_r21_c2;
    wire stage0_r22_c1;
    wire stage0_r23_c0;
    wire stage0_r0_c24;
    wire stage0_r1_c23;
    wire stage0_r2_c22;
    wire stage0_r3_c21;
    wire stage0_r4_c20;
    wire stage0_r5_c19;
    wire stage0_r6_c18;
    wire stage0_r7_c17;
    wire stage0_r8_c16;
    wire stage0_r9_c15;
    wire stage0_r10_c14;
    wire stage0_r11_c13;
    wire stage0_r12_c12;
    wire stage0_r13_c11;
    wire stage0_r14_c10;
    wire stage0_r15_c9;
    wire stage0_r16_c8;
    wire stage0_r17_c7;
    wire stage0_r18_c6;
    wire stage0_r19_c5;
    wire stage0_r20_c4;
    wire stage0_r21_c3;
    wire stage0_r22_c2;
    wire stage0_r23_c1;
    wire stage0_r24_c0;
    wire stage0_r0_c25;
    wire stage0_r1_c24;
    wire stage0_r2_c23;
    wire stage0_r3_c22;
    wire stage0_r4_c21;
    wire stage0_r5_c20;
    wire stage0_r6_c19;
    wire stage0_r7_c18;
    wire stage0_r8_c17;
    wire stage0_r9_c16;
    wire stage0_r10_c15;
    wire stage0_r11_c14;
    wire stage0_r12_c13;
    wire stage0_r13_c12;
    wire stage0_r14_c11;
    wire stage0_r15_c10;
    wire stage0_r16_c9;
    wire stage0_r17_c8;
    wire stage0_r18_c7;
    wire stage0_r19_c6;
    wire stage0_r20_c5;
    wire stage0_r21_c4;
    wire stage0_r22_c3;
    wire stage0_r23_c2;
    wire stage0_r24_c1;
    wire stage0_r25_c0;
    wire stage0_r0_c26;
    wire stage0_r1_c25;
    wire stage0_r2_c24;
    wire stage0_r3_c23;
    wire stage0_r4_c22;
    wire stage0_r5_c21;
    wire stage0_r6_c20;
    wire stage0_r7_c19;
    wire stage0_r8_c18;
    wire stage0_r9_c17;
    wire stage0_r10_c16;
    wire stage0_r11_c15;
    wire stage0_r12_c14;
    wire stage0_r13_c13;
    wire stage0_r14_c12;
    wire stage0_r15_c11;
    wire stage0_r16_c10;
    wire stage0_r17_c9;
    wire stage0_r18_c8;
    wire stage0_r19_c7;
    wire stage0_r20_c6;
    wire stage0_r21_c5;
    wire stage0_r22_c4;
    wire stage0_r23_c3;
    wire stage0_r24_c2;
    wire stage0_r25_c1;
    wire stage0_r26_c0;
    wire stage0_r0_c27;
    wire stage0_r1_c26;
    wire stage0_r2_c25;
    wire stage0_r3_c24;
    wire stage0_r4_c23;
    wire stage0_r5_c22;
    wire stage0_r6_c21;
    wire stage0_r7_c20;
    wire stage0_r8_c19;
    wire stage0_r9_c18;
    wire stage0_r10_c17;
    wire stage0_r11_c16;
    wire stage0_r12_c15;
    wire stage0_r13_c14;
    wire stage0_r14_c13;
    wire stage0_r15_c12;
    wire stage0_r16_c11;
    wire stage0_r17_c10;
    wire stage0_r18_c9;
    wire stage0_r19_c8;
    wire stage0_r20_c7;
    wire stage0_r21_c6;
    wire stage0_r22_c5;
    wire stage0_r23_c4;
    wire stage0_r24_c3;
    wire stage0_r25_c2;
    wire stage0_r26_c1;
    wire stage0_r27_c0;
    wire stage0_r0_c28;
    wire stage0_r1_c27;
    wire stage0_r2_c26;
    wire stage0_r3_c25;
    wire stage0_r4_c24;
    wire stage0_r5_c23;
    wire stage0_r6_c22;
    wire stage0_r7_c21;
    wire stage0_r8_c20;
    wire stage0_r9_c19;
    wire stage0_r10_c18;
    wire stage0_r11_c17;
    wire stage0_r12_c16;
    wire stage0_r13_c15;
    wire stage0_r14_c14;
    wire stage0_r15_c13;
    wire stage0_r16_c12;
    wire stage0_r17_c11;
    wire stage0_r18_c10;
    wire stage0_r19_c9;
    wire stage0_r20_c8;
    wire stage0_r21_c7;
    wire stage0_r22_c6;
    wire stage0_r23_c5;
    wire stage0_r24_c4;
    wire stage0_r25_c3;
    wire stage0_r26_c2;
    wire stage0_r27_c1;
    wire stage0_r28_c0;
    wire stage0_r0_c29;
    wire stage0_r1_c28;
    wire stage0_r2_c27;
    wire stage0_r3_c26;
    wire stage0_r4_c25;
    wire stage0_r5_c24;
    wire stage0_r6_c23;
    wire stage0_r7_c22;
    wire stage0_r8_c21;
    wire stage0_r9_c20;
    wire stage0_r10_c19;
    wire stage0_r11_c18;
    wire stage0_r12_c17;
    wire stage0_r13_c16;
    wire stage0_r14_c15;
    wire stage0_r15_c14;
    wire stage0_r16_c13;
    wire stage0_r17_c12;
    wire stage0_r18_c11;
    wire stage0_r19_c10;
    wire stage0_r20_c9;
    wire stage0_r21_c8;
    wire stage0_r22_c7;
    wire stage0_r23_c6;
    wire stage0_r24_c5;
    wire stage0_r25_c4;
    wire stage0_r26_c3;
    wire stage0_r27_c2;
    wire stage0_r28_c1;
    wire stage0_r29_c0;
    wire stage0_r0_c30;
    wire stage0_r1_c29;
    wire stage0_r2_c28;
    wire stage0_r3_c27;
    wire stage0_r4_c26;
    wire stage0_r5_c25;
    wire stage0_r6_c24;
    wire stage0_r7_c23;
    wire stage0_r8_c22;
    wire stage0_r9_c21;
    wire stage0_r10_c20;
    wire stage0_r11_c19;
    wire stage0_r12_c18;
    wire stage0_r13_c17;
    wire stage0_r14_c16;
    wire stage0_r15_c15;
    wire stage0_r16_c14;
    wire stage0_r17_c13;
    wire stage0_r18_c12;
    wire stage0_r19_c11;
    wire stage0_r20_c10;
    wire stage0_r21_c9;
    wire stage0_r22_c8;
    wire stage0_r23_c7;
    wire stage0_r24_c6;
    wire stage0_r25_c5;
    wire stage0_r26_c4;
    wire stage0_r27_c3;
    wire stage0_r28_c2;
    wire stage0_r29_c1;
    wire stage0_r30_c0;
    wire stage0_r0_c31;
    wire stage0_r1_c30;
    wire stage0_r2_c29;
    wire stage0_r3_c28;
    wire stage0_r4_c27;
    wire stage0_r5_c26;
    wire stage0_r6_c25;
    wire stage0_r7_c24;
    wire stage0_r8_c23;
    wire stage0_r9_c22;
    wire stage0_r10_c21;
    wire stage0_r11_c20;
    wire stage0_r12_c19;
    wire stage0_r13_c18;
    wire stage0_r14_c17;
    wire stage0_r15_c16;
    wire stage0_r16_c15;
    wire stage0_r17_c14;
    wire stage0_r18_c13;
    wire stage0_r19_c12;
    wire stage0_r20_c11;
    wire stage0_r21_c10;
    wire stage0_r22_c9;
    wire stage0_r23_c8;
    wire stage0_r24_c7;
    wire stage0_r25_c6;
    wire stage0_r26_c5;
    wire stage0_r27_c4;
    wire stage0_r28_c3;
    wire stage0_r29_c2;
    wire stage0_r30_c1;
    wire stage0_r31_c0;
    wire stage0_r0_c32;
    wire stage0_r1_c31;
    wire stage0_r2_c30;
    wire stage0_r3_c29;
    wire stage0_r4_c28;
    wire stage0_r5_c27;
    wire stage0_r6_c26;
    wire stage0_r7_c25;
    wire stage0_r8_c24;
    wire stage0_r9_c23;
    wire stage0_r10_c22;
    wire stage0_r11_c21;
    wire stage0_r12_c20;
    wire stage0_r13_c19;
    wire stage0_r14_c18;
    wire stage0_r15_c17;
    wire stage0_r16_c16;
    wire stage0_r17_c15;
    wire stage0_r18_c14;
    wire stage0_r19_c13;
    wire stage0_r20_c12;
    wire stage0_r21_c11;
    wire stage0_r22_c10;
    wire stage0_r23_c9;
    wire stage0_r24_c8;
    wire stage0_r25_c7;
    wire stage0_r26_c6;
    wire stage0_r27_c5;
    wire stage0_r28_c4;
    wire stage0_r29_c3;
    wire stage0_r30_c2;
    wire stage0_r31_c1;
    wire stage0_r32_c0;
    wire stage0_r0_c33;
    wire stage0_r1_c32;
    wire stage0_r2_c31;
    wire stage0_r3_c30;
    wire stage0_r4_c29;
    wire stage0_r5_c28;
    wire stage0_r6_c27;
    wire stage0_r7_c26;
    wire stage0_r8_c25;
    wire stage0_r9_c24;
    wire stage0_r10_c23;
    wire stage0_r11_c22;
    wire stage0_r12_c21;
    wire stage0_r13_c20;
    wire stage0_r14_c19;
    wire stage0_r15_c18;
    wire stage0_r16_c17;
    wire stage0_r17_c16;
    wire stage0_r18_c15;
    wire stage0_r19_c14;
    wire stage0_r20_c13;
    wire stage0_r21_c12;
    wire stage0_r22_c11;
    wire stage0_r23_c10;
    wire stage0_r24_c9;
    wire stage0_r25_c8;
    wire stage0_r26_c7;
    wire stage0_r27_c6;
    wire stage0_r28_c5;
    wire stage0_r29_c4;
    wire stage0_r30_c3;
    wire stage0_r31_c2;
    wire stage0_r32_c1;
    wire stage0_r33_c0;
    wire stage0_r0_c34;
    wire stage0_r1_c33;
    wire stage0_r2_c32;
    wire stage0_r3_c31;
    wire stage0_r4_c30;
    wire stage0_r5_c29;
    wire stage0_r6_c28;
    wire stage0_r7_c27;
    wire stage0_r8_c26;
    wire stage0_r9_c25;
    wire stage0_r10_c24;
    wire stage0_r11_c23;
    wire stage0_r12_c22;
    wire stage0_r13_c21;
    wire stage0_r14_c20;
    wire stage0_r15_c19;
    wire stage0_r16_c18;
    wire stage0_r17_c17;
    wire stage0_r18_c16;
    wire stage0_r19_c15;
    wire stage0_r20_c14;
    wire stage0_r21_c13;
    wire stage0_r22_c12;
    wire stage0_r23_c11;
    wire stage0_r24_c10;
    wire stage0_r25_c9;
    wire stage0_r26_c8;
    wire stage0_r27_c7;
    wire stage0_r28_c6;
    wire stage0_r29_c5;
    wire stage0_r30_c4;
    wire stage0_r31_c3;
    wire stage0_r32_c2;
    wire stage0_r33_c1;
    wire stage0_r34_c0;
    wire stage0_r0_c35;
    wire stage0_r1_c34;
    wire stage0_r2_c33;
    wire stage0_r3_c32;
    wire stage0_r4_c31;
    wire stage0_r5_c30;
    wire stage0_r6_c29;
    wire stage0_r7_c28;
    wire stage0_r8_c27;
    wire stage0_r9_c26;
    wire stage0_r10_c25;
    wire stage0_r11_c24;
    wire stage0_r12_c23;
    wire stage0_r13_c22;
    wire stage0_r14_c21;
    wire stage0_r15_c20;
    wire stage0_r16_c19;
    wire stage0_r17_c18;
    wire stage0_r18_c17;
    wire stage0_r19_c16;
    wire stage0_r20_c15;
    wire stage0_r21_c14;
    wire stage0_r22_c13;
    wire stage0_r23_c12;
    wire stage0_r24_c11;
    wire stage0_r25_c10;
    wire stage0_r26_c9;
    wire stage0_r27_c8;
    wire stage0_r28_c7;
    wire stage0_r29_c6;
    wire stage0_r30_c5;
    wire stage0_r31_c4;
    wire stage0_r32_c3;
    wire stage0_r33_c2;
    wire stage0_r34_c1;
    wire stage0_r35_c0;
    wire stage0_r0_c36;
    wire stage0_r1_c35;
    wire stage0_r2_c34;
    wire stage0_r3_c33;
    wire stage0_r4_c32;
    wire stage0_r5_c31;
    wire stage0_r6_c30;
    wire stage0_r7_c29;
    wire stage0_r8_c28;
    wire stage0_r9_c27;
    wire stage0_r10_c26;
    wire stage0_r11_c25;
    wire stage0_r12_c24;
    wire stage0_r13_c23;
    wire stage0_r14_c22;
    wire stage0_r15_c21;
    wire stage0_r16_c20;
    wire stage0_r17_c19;
    wire stage0_r18_c18;
    wire stage0_r19_c17;
    wire stage0_r20_c16;
    wire stage0_r21_c15;
    wire stage0_r22_c14;
    wire stage0_r23_c13;
    wire stage0_r24_c12;
    wire stage0_r25_c11;
    wire stage0_r26_c10;
    wire stage0_r27_c9;
    wire stage0_r28_c8;
    wire stage0_r29_c7;
    wire stage0_r30_c6;
    wire stage0_r31_c5;
    wire stage0_r32_c4;
    wire stage0_r33_c3;
    wire stage0_r34_c2;
    wire stage0_r35_c1;
    wire stage0_r36_c0;
    wire stage0_r0_c37;
    wire stage0_r1_c36;
    wire stage0_r2_c35;
    wire stage0_r3_c34;
    wire stage0_r4_c33;
    wire stage0_r5_c32;
    wire stage0_r6_c31;
    wire stage0_r7_c30;
    wire stage0_r8_c29;
    wire stage0_r9_c28;
    wire stage0_r10_c27;
    wire stage0_r11_c26;
    wire stage0_r12_c25;
    wire stage0_r13_c24;
    wire stage0_r14_c23;
    wire stage0_r15_c22;
    wire stage0_r16_c21;
    wire stage0_r17_c20;
    wire stage0_r18_c19;
    wire stage0_r19_c18;
    wire stage0_r20_c17;
    wire stage0_r21_c16;
    wire stage0_r22_c15;
    wire stage0_r23_c14;
    wire stage0_r24_c13;
    wire stage0_r25_c12;
    wire stage0_r26_c11;
    wire stage0_r27_c10;
    wire stage0_r28_c9;
    wire stage0_r29_c8;
    wire stage0_r30_c7;
    wire stage0_r31_c6;
    wire stage0_r32_c5;
    wire stage0_r33_c4;
    wire stage0_r34_c3;
    wire stage0_r35_c2;
    wire stage0_r36_c1;
    wire stage0_r37_c0;
    wire stage0_r0_c38;
    wire stage0_r1_c37;
    wire stage0_r2_c36;
    wire stage0_r3_c35;
    wire stage0_r4_c34;
    wire stage0_r5_c33;
    wire stage0_r6_c32;
    wire stage0_r7_c31;
    wire stage0_r8_c30;
    wire stage0_r9_c29;
    wire stage0_r10_c28;
    wire stage0_r11_c27;
    wire stage0_r12_c26;
    wire stage0_r13_c25;
    wire stage0_r14_c24;
    wire stage0_r15_c23;
    wire stage0_r16_c22;
    wire stage0_r17_c21;
    wire stage0_r18_c20;
    wire stage0_r19_c19;
    wire stage0_r20_c18;
    wire stage0_r21_c17;
    wire stage0_r22_c16;
    wire stage0_r23_c15;
    wire stage0_r24_c14;
    wire stage0_r25_c13;
    wire stage0_r26_c12;
    wire stage0_r27_c11;
    wire stage0_r28_c10;
    wire stage0_r29_c9;
    wire stage0_r30_c8;
    wire stage0_r31_c7;
    wire stage0_r32_c6;
    wire stage0_r33_c5;
    wire stage0_r34_c4;
    wire stage0_r35_c3;
    wire stage0_r36_c2;
    wire stage0_r37_c1;
    wire stage0_r38_c0;
    wire stage0_r0_c39;
    wire stage0_r1_c38;
    wire stage0_r2_c37;
    wire stage0_r3_c36;
    wire stage0_r4_c35;
    wire stage0_r5_c34;
    wire stage0_r6_c33;
    wire stage0_r7_c32;
    wire stage0_r8_c31;
    wire stage0_r9_c30;
    wire stage0_r10_c29;
    wire stage0_r11_c28;
    wire stage0_r12_c27;
    wire stage0_r13_c26;
    wire stage0_r14_c25;
    wire stage0_r15_c24;
    wire stage0_r16_c23;
    wire stage0_r17_c22;
    wire stage0_r18_c21;
    wire stage0_r19_c20;
    wire stage0_r20_c19;
    wire stage0_r21_c18;
    wire stage0_r22_c17;
    wire stage0_r23_c16;
    wire stage0_r24_c15;
    wire stage0_r25_c14;
    wire stage0_r26_c13;
    wire stage0_r27_c12;
    wire stage0_r28_c11;
    wire stage0_r29_c10;
    wire stage0_r30_c9;
    wire stage0_r31_c8;
    wire stage0_r32_c7;
    wire stage0_r33_c6;
    wire stage0_r34_c5;
    wire stage0_r35_c4;
    wire stage0_r36_c3;
    wire stage0_r37_c2;
    wire stage0_r38_c1;
    wire stage0_r39_c0;
    wire stage0_r0_c40;
    wire stage0_r1_c39;
    wire stage0_r2_c38;
    wire stage0_r3_c37;
    wire stage0_r4_c36;
    wire stage0_r5_c35;
    wire stage0_r6_c34;
    wire stage0_r7_c33;
    wire stage0_r8_c32;
    wire stage0_r9_c31;
    wire stage0_r10_c30;
    wire stage0_r11_c29;
    wire stage0_r12_c28;
    wire stage0_r13_c27;
    wire stage0_r14_c26;
    wire stage0_r15_c25;
    wire stage0_r16_c24;
    wire stage0_r17_c23;
    wire stage0_r18_c22;
    wire stage0_r19_c21;
    wire stage0_r20_c20;
    wire stage0_r21_c19;
    wire stage0_r22_c18;
    wire stage0_r23_c17;
    wire stage0_r24_c16;
    wire stage0_r25_c15;
    wire stage0_r26_c14;
    wire stage0_r27_c13;
    wire stage0_r28_c12;
    wire stage0_r29_c11;
    wire stage0_r30_c10;
    wire stage0_r31_c9;
    wire stage0_r32_c8;
    wire stage0_r33_c7;
    wire stage0_r34_c6;
    wire stage0_r35_c5;
    wire stage0_r36_c4;
    wire stage0_r37_c3;
    wire stage0_r38_c2;
    wire stage0_r39_c1;
    wire stage0_r40_c0;
    wire stage0_r1_c40;
    wire stage0_r2_c39;
    wire stage0_r3_c38;
    wire stage0_r4_c37;
    wire stage0_r5_c36;
    wire stage0_r6_c35;
    wire stage0_r7_c34;
    wire stage0_r8_c33;
    wire stage0_r9_c32;
    wire stage0_r10_c31;
    wire stage0_r11_c30;
    wire stage0_r12_c29;
    wire stage0_r13_c28;
    wire stage0_r14_c27;
    wire stage0_r15_c26;
    wire stage0_r16_c25;
    wire stage0_r17_c24;
    wire stage0_r18_c23;
    wire stage0_r19_c22;
    wire stage0_r20_c21;
    wire stage0_r21_c20;
    wire stage0_r22_c19;
    wire stage0_r23_c18;
    wire stage0_r24_c17;
    wire stage0_r25_c16;
    wire stage0_r26_c15;
    wire stage0_r27_c14;
    wire stage0_r28_c13;
    wire stage0_r29_c12;
    wire stage0_r30_c11;
    wire stage0_r31_c10;
    wire stage0_r32_c9;
    wire stage0_r33_c8;
    wire stage0_r34_c7;
    wire stage0_r35_c6;
    wire stage0_r36_c5;
    wire stage0_r37_c4;
    wire stage0_r38_c3;
    wire stage0_r39_c2;
    wire stage0_r40_c1;
    wire stage0_r41_c0;
    wire stage0_r2_c40;
    wire stage0_r3_c39;
    wire stage0_r4_c38;
    wire stage0_r5_c37;
    wire stage0_r6_c36;
    wire stage0_r7_c35;
    wire stage0_r8_c34;
    wire stage0_r9_c33;
    wire stage0_r10_c32;
    wire stage0_r11_c31;
    wire stage0_r12_c30;
    wire stage0_r13_c29;
    wire stage0_r14_c28;
    wire stage0_r15_c27;
    wire stage0_r16_c26;
    wire stage0_r17_c25;
    wire stage0_r18_c24;
    wire stage0_r19_c23;
    wire stage0_r20_c22;
    wire stage0_r21_c21;
    wire stage0_r22_c20;
    wire stage0_r23_c19;
    wire stage0_r24_c18;
    wire stage0_r25_c17;
    wire stage0_r26_c16;
    wire stage0_r27_c15;
    wire stage0_r28_c14;
    wire stage0_r29_c13;
    wire stage0_r30_c12;
    wire stage0_r31_c11;
    wire stage0_r32_c10;
    wire stage0_r33_c9;
    wire stage0_r34_c8;
    wire stage0_r35_c7;
    wire stage0_r36_c6;
    wire stage0_r37_c5;
    wire stage0_r38_c4;
    wire stage0_r39_c3;
    wire stage0_r40_c2;
    wire stage0_r41_c1;
    wire stage0_r42_c0;
    wire stage0_r3_c40;
    wire stage0_r4_c39;
    wire stage0_r5_c38;
    wire stage0_r6_c37;
    wire stage0_r7_c36;
    wire stage0_r8_c35;
    wire stage0_r9_c34;
    wire stage0_r10_c33;
    wire stage0_r11_c32;
    wire stage0_r12_c31;
    wire stage0_r13_c30;
    wire stage0_r14_c29;
    wire stage0_r15_c28;
    wire stage0_r16_c27;
    wire stage0_r17_c26;
    wire stage0_r18_c25;
    wire stage0_r19_c24;
    wire stage0_r20_c23;
    wire stage0_r21_c22;
    wire stage0_r22_c21;
    wire stage0_r23_c20;
    wire stage0_r24_c19;
    wire stage0_r25_c18;
    wire stage0_r26_c17;
    wire stage0_r27_c16;
    wire stage0_r28_c15;
    wire stage0_r29_c14;
    wire stage0_r30_c13;
    wire stage0_r31_c12;
    wire stage0_r32_c11;
    wire stage0_r33_c10;
    wire stage0_r34_c9;
    wire stage0_r35_c8;
    wire stage0_r36_c7;
    wire stage0_r37_c6;
    wire stage0_r38_c5;
    wire stage0_r39_c4;
    wire stage0_r40_c3;
    wire stage0_r41_c2;
    wire stage0_r42_c1;
    wire stage0_r43_c0;
    wire stage0_r4_c40;
    wire stage0_r5_c39;
    wire stage0_r6_c38;
    wire stage0_r7_c37;
    wire stage0_r8_c36;
    wire stage0_r9_c35;
    wire stage0_r10_c34;
    wire stage0_r11_c33;
    wire stage0_r12_c32;
    wire stage0_r13_c31;
    wire stage0_r14_c30;
    wire stage0_r15_c29;
    wire stage0_r16_c28;
    wire stage0_r17_c27;
    wire stage0_r18_c26;
    wire stage0_r19_c25;
    wire stage0_r20_c24;
    wire stage0_r21_c23;
    wire stage0_r22_c22;
    wire stage0_r23_c21;
    wire stage0_r24_c20;
    wire stage0_r25_c19;
    wire stage0_r26_c18;
    wire stage0_r27_c17;
    wire stage0_r28_c16;
    wire stage0_r29_c15;
    wire stage0_r30_c14;
    wire stage0_r31_c13;
    wire stage0_r32_c12;
    wire stage0_r33_c11;
    wire stage0_r34_c10;
    wire stage0_r35_c9;
    wire stage0_r36_c8;
    wire stage0_r37_c7;
    wire stage0_r38_c6;
    wire stage0_r39_c5;
    wire stage0_r40_c4;
    wire stage0_r41_c3;
    wire stage0_r42_c2;
    wire stage0_r43_c1;
    wire stage0_r44_c0;
    wire stage0_r5_c40;
    wire stage0_r6_c39;
    wire stage0_r7_c38;
    wire stage0_r8_c37;
    wire stage0_r9_c36;
    wire stage0_r10_c35;
    wire stage0_r11_c34;
    wire stage0_r12_c33;
    wire stage0_r13_c32;
    wire stage0_r14_c31;
    wire stage0_r15_c30;
    wire stage0_r16_c29;
    wire stage0_r17_c28;
    wire stage0_r18_c27;
    wire stage0_r19_c26;
    wire stage0_r20_c25;
    wire stage0_r21_c24;
    wire stage0_r22_c23;
    wire stage0_r23_c22;
    wire stage0_r24_c21;
    wire stage0_r25_c20;
    wire stage0_r26_c19;
    wire stage0_r27_c18;
    wire stage0_r28_c17;
    wire stage0_r29_c16;
    wire stage0_r30_c15;
    wire stage0_r31_c14;
    wire stage0_r32_c13;
    wire stage0_r33_c12;
    wire stage0_r34_c11;
    wire stage0_r35_c10;
    wire stage0_r36_c9;
    wire stage0_r37_c8;
    wire stage0_r38_c7;
    wire stage0_r39_c6;
    wire stage0_r40_c5;
    wire stage0_r41_c4;
    wire stage0_r42_c3;
    wire stage0_r43_c2;
    wire stage0_r44_c1;
    wire stage0_r45_c0;
    wire stage0_r6_c40;
    wire stage0_r7_c39;
    wire stage0_r8_c38;
    wire stage0_r9_c37;
    wire stage0_r10_c36;
    wire stage0_r11_c35;
    wire stage0_r12_c34;
    wire stage0_r13_c33;
    wire stage0_r14_c32;
    wire stage0_r15_c31;
    wire stage0_r16_c30;
    wire stage0_r17_c29;
    wire stage0_r18_c28;
    wire stage0_r19_c27;
    wire stage0_r20_c26;
    wire stage0_r21_c25;
    wire stage0_r22_c24;
    wire stage0_r23_c23;
    wire stage0_r24_c22;
    wire stage0_r25_c21;
    wire stage0_r26_c20;
    wire stage0_r27_c19;
    wire stage0_r28_c18;
    wire stage0_r29_c17;
    wire stage0_r30_c16;
    wire stage0_r31_c15;
    wire stage0_r32_c14;
    wire stage0_r33_c13;
    wire stage0_r34_c12;
    wire stage0_r35_c11;
    wire stage0_r36_c10;
    wire stage0_r37_c9;
    wire stage0_r38_c8;
    wire stage0_r39_c7;
    wire stage0_r40_c6;
    wire stage0_r41_c5;
    wire stage0_r42_c4;
    wire stage0_r43_c3;
    wire stage0_r44_c2;
    wire stage0_r45_c1;
    wire stage0_r46_c0;
    wire stage0_r7_c40;
    wire stage0_r8_c39;
    wire stage0_r9_c38;
    wire stage0_r10_c37;
    wire stage0_r11_c36;
    wire stage0_r12_c35;
    wire stage0_r13_c34;
    wire stage0_r14_c33;
    wire stage0_r15_c32;
    wire stage0_r16_c31;
    wire stage0_r17_c30;
    wire stage0_r18_c29;
    wire stage0_r19_c28;
    wire stage0_r20_c27;
    wire stage0_r21_c26;
    wire stage0_r22_c25;
    wire stage0_r23_c24;
    wire stage0_r24_c23;
    wire stage0_r25_c22;
    wire stage0_r26_c21;
    wire stage0_r27_c20;
    wire stage0_r28_c19;
    wire stage0_r29_c18;
    wire stage0_r30_c17;
    wire stage0_r31_c16;
    wire stage0_r32_c15;
    wire stage0_r33_c14;
    wire stage0_r34_c13;
    wire stage0_r35_c12;
    wire stage0_r36_c11;
    wire stage0_r37_c10;
    wire stage0_r38_c9;
    wire stage0_r39_c8;
    wire stage0_r40_c7;
    wire stage0_r41_c6;
    wire stage0_r42_c5;
    wire stage0_r43_c4;
    wire stage0_r44_c3;
    wire stage0_r45_c2;
    wire stage0_r46_c1;
    wire stage0_r47_c0;
    wire stage0_r8_c40;
    wire stage0_r9_c39;
    wire stage0_r10_c38;
    wire stage0_r11_c37;
    wire stage0_r12_c36;
    wire stage0_r13_c35;
    wire stage0_r14_c34;
    wire stage0_r15_c33;
    wire stage0_r16_c32;
    wire stage0_r17_c31;
    wire stage0_r18_c30;
    wire stage0_r19_c29;
    wire stage0_r20_c28;
    wire stage0_r21_c27;
    wire stage0_r22_c26;
    wire stage0_r23_c25;
    wire stage0_r24_c24;
    wire stage0_r25_c23;
    wire stage0_r26_c22;
    wire stage0_r27_c21;
    wire stage0_r28_c20;
    wire stage0_r29_c19;
    wire stage0_r30_c18;
    wire stage0_r31_c17;
    wire stage0_r32_c16;
    wire stage0_r33_c15;
    wire stage0_r34_c14;
    wire stage0_r35_c13;
    wire stage0_r36_c12;
    wire stage0_r37_c11;
    wire stage0_r38_c10;
    wire stage0_r39_c9;
    wire stage0_r40_c8;
    wire stage0_r41_c7;
    wire stage0_r42_c6;
    wire stage0_r43_c5;
    wire stage0_r44_c4;
    wire stage0_r45_c3;
    wire stage0_r46_c2;
    wire stage0_r47_c1;
    wire stage0_r48_c0;
    wire stage0_r9_c40;
    wire stage0_r10_c39;
    wire stage0_r11_c38;
    wire stage0_r12_c37;
    wire stage0_r13_c36;
    wire stage0_r14_c35;
    wire stage0_r15_c34;
    wire stage0_r16_c33;
    wire stage0_r17_c32;
    wire stage0_r18_c31;
    wire stage0_r19_c30;
    wire stage0_r20_c29;
    wire stage0_r21_c28;
    wire stage0_r22_c27;
    wire stage0_r23_c26;
    wire stage0_r24_c25;
    wire stage0_r25_c24;
    wire stage0_r26_c23;
    wire stage0_r27_c22;
    wire stage0_r28_c21;
    wire stage0_r29_c20;
    wire stage0_r30_c19;
    wire stage0_r31_c18;
    wire stage0_r32_c17;
    wire stage0_r33_c16;
    wire stage0_r34_c15;
    wire stage0_r35_c14;
    wire stage0_r36_c13;
    wire stage0_r37_c12;
    wire stage0_r38_c11;
    wire stage0_r39_c10;
    wire stage0_r40_c9;
    wire stage0_r41_c8;
    wire stage0_r42_c7;
    wire stage0_r43_c6;
    wire stage0_r44_c5;
    wire stage0_r45_c4;
    wire stage0_r46_c3;
    wire stage0_r47_c2;
    wire stage0_r48_c1;
    wire stage0_r49_c0;
    wire stage0_r10_c40;
    wire stage0_r11_c39;
    wire stage0_r12_c38;
    wire stage0_r13_c37;
    wire stage0_r14_c36;
    wire stage0_r15_c35;
    wire stage0_r16_c34;
    wire stage0_r17_c33;
    wire stage0_r18_c32;
    wire stage0_r19_c31;
    wire stage0_r20_c30;
    wire stage0_r21_c29;
    wire stage0_r22_c28;
    wire stage0_r23_c27;
    wire stage0_r24_c26;
    wire stage0_r25_c25;
    wire stage0_r26_c24;
    wire stage0_r27_c23;
    wire stage0_r28_c22;
    wire stage0_r29_c21;
    wire stage0_r30_c20;
    wire stage0_r31_c19;
    wire stage0_r32_c18;
    wire stage0_r33_c17;
    wire stage0_r34_c16;
    wire stage0_r35_c15;
    wire stage0_r36_c14;
    wire stage0_r37_c13;
    wire stage0_r38_c12;
    wire stage0_r39_c11;
    wire stage0_r40_c10;
    wire stage0_r41_c9;
    wire stage0_r42_c8;
    wire stage0_r43_c7;
    wire stage0_r44_c6;
    wire stage0_r45_c5;
    wire stage0_r46_c4;
    wire stage0_r47_c3;
    wire stage0_r48_c2;
    wire stage0_r49_c1;
    wire stage0_r50_c0;
    wire stage0_r11_c40;
    wire stage0_r12_c39;
    wire stage0_r13_c38;
    wire stage0_r14_c37;
    wire stage0_r15_c36;
    wire stage0_r16_c35;
    wire stage0_r17_c34;
    wire stage0_r18_c33;
    wire stage0_r19_c32;
    wire stage0_r20_c31;
    wire stage0_r21_c30;
    wire stage0_r22_c29;
    wire stage0_r23_c28;
    wire stage0_r24_c27;
    wire stage0_r25_c26;
    wire stage0_r26_c25;
    wire stage0_r27_c24;
    wire stage0_r28_c23;
    wire stage0_r29_c22;
    wire stage0_r30_c21;
    wire stage0_r31_c20;
    wire stage0_r32_c19;
    wire stage0_r33_c18;
    wire stage0_r34_c17;
    wire stage0_r35_c16;
    wire stage0_r36_c15;
    wire stage0_r37_c14;
    wire stage0_r38_c13;
    wire stage0_r39_c12;
    wire stage0_r40_c11;
    wire stage0_r41_c10;
    wire stage0_r42_c9;
    wire stage0_r43_c8;
    wire stage0_r44_c7;
    wire stage0_r45_c6;
    wire stage0_r46_c5;
    wire stage0_r47_c4;
    wire stage0_r48_c3;
    wire stage0_r49_c2;
    wire stage0_r50_c1;
    wire stage0_r51_c0;
    wire stage0_r12_c40;
    wire stage0_r13_c39;
    wire stage0_r14_c38;
    wire stage0_r15_c37;
    wire stage0_r16_c36;
    wire stage0_r17_c35;
    wire stage0_r18_c34;
    wire stage0_r19_c33;
    wire stage0_r20_c32;
    wire stage0_r21_c31;
    wire stage0_r22_c30;
    wire stage0_r23_c29;
    wire stage0_r24_c28;
    wire stage0_r25_c27;
    wire stage0_r26_c26;
    wire stage0_r27_c25;
    wire stage0_r28_c24;
    wire stage0_r29_c23;
    wire stage0_r30_c22;
    wire stage0_r31_c21;
    wire stage0_r32_c20;
    wire stage0_r33_c19;
    wire stage0_r34_c18;
    wire stage0_r35_c17;
    wire stage0_r36_c16;
    wire stage0_r37_c15;
    wire stage0_r38_c14;
    wire stage0_r39_c13;
    wire stage0_r40_c12;
    wire stage0_r41_c11;
    wire stage0_r42_c10;
    wire stage0_r43_c9;
    wire stage0_r44_c8;
    wire stage0_r45_c7;
    wire stage0_r46_c6;
    wire stage0_r47_c5;
    wire stage0_r48_c4;
    wire stage0_r49_c3;
    wire stage0_r50_c2;
    wire stage0_r51_c1;
    wire stage0_r52_c0;
    wire stage0_r13_c40;
    wire stage0_r14_c39;
    wire stage0_r15_c38;
    wire stage0_r16_c37;
    wire stage0_r17_c36;
    wire stage0_r18_c35;
    wire stage0_r19_c34;
    wire stage0_r20_c33;
    wire stage0_r21_c32;
    wire stage0_r22_c31;
    wire stage0_r23_c30;
    wire stage0_r24_c29;
    wire stage0_r25_c28;
    wire stage0_r26_c27;
    wire stage0_r27_c26;
    wire stage0_r28_c25;
    wire stage0_r29_c24;
    wire stage0_r30_c23;
    wire stage0_r31_c22;
    wire stage0_r32_c21;
    wire stage0_r33_c20;
    wire stage0_r34_c19;
    wire stage0_r35_c18;
    wire stage0_r36_c17;
    wire stage0_r37_c16;
    wire stage0_r38_c15;
    wire stage0_r39_c14;
    wire stage0_r40_c13;
    wire stage0_r41_c12;
    wire stage0_r42_c11;
    wire stage0_r43_c10;
    wire stage0_r44_c9;
    wire stage0_r45_c8;
    wire stage0_r46_c7;
    wire stage0_r47_c6;
    wire stage0_r48_c5;
    wire stage0_r49_c4;
    wire stage0_r50_c3;
    wire stage0_r51_c2;
    wire stage0_r52_c1;
    wire stage0_r53_c0;
    wire stage0_r14_c40;
    wire stage0_r15_c39;
    wire stage0_r16_c38;
    wire stage0_r17_c37;
    wire stage0_r18_c36;
    wire stage0_r19_c35;
    wire stage0_r20_c34;
    wire stage0_r21_c33;
    wire stage0_r22_c32;
    wire stage0_r23_c31;
    wire stage0_r24_c30;
    wire stage0_r25_c29;
    wire stage0_r26_c28;
    wire stage0_r27_c27;
    wire stage0_r28_c26;
    wire stage0_r29_c25;
    wire stage0_r30_c24;
    wire stage0_r31_c23;
    wire stage0_r32_c22;
    wire stage0_r33_c21;
    wire stage0_r34_c20;
    wire stage0_r35_c19;
    wire stage0_r36_c18;
    wire stage0_r37_c17;
    wire stage0_r38_c16;
    wire stage0_r39_c15;
    wire stage0_r40_c14;
    wire stage0_r41_c13;
    wire stage0_r42_c12;
    wire stage0_r43_c11;
    wire stage0_r44_c10;
    wire stage0_r45_c9;
    wire stage0_r46_c8;
    wire stage0_r47_c7;
    wire stage0_r48_c6;
    wire stage0_r49_c5;
    wire stage0_r50_c4;
    wire stage0_r51_c3;
    wire stage0_r52_c2;
    wire stage0_r53_c1;
    wire stage0_r54_c0;
    wire stage0_r15_c40;
    wire stage0_r16_c39;
    wire stage0_r17_c38;
    wire stage0_r18_c37;
    wire stage0_r19_c36;
    wire stage0_r20_c35;
    wire stage0_r21_c34;
    wire stage0_r22_c33;
    wire stage0_r23_c32;
    wire stage0_r24_c31;
    wire stage0_r25_c30;
    wire stage0_r26_c29;
    wire stage0_r27_c28;
    wire stage0_r28_c27;
    wire stage0_r29_c26;
    wire stage0_r30_c25;
    wire stage0_r31_c24;
    wire stage0_r32_c23;
    wire stage0_r33_c22;
    wire stage0_r34_c21;
    wire stage0_r35_c20;
    wire stage0_r36_c19;
    wire stage0_r37_c18;
    wire stage0_r38_c17;
    wire stage0_r39_c16;
    wire stage0_r40_c15;
    wire stage0_r41_c14;
    wire stage0_r42_c13;
    wire stage0_r43_c12;
    wire stage0_r44_c11;
    wire stage0_r45_c10;
    wire stage0_r46_c9;
    wire stage0_r47_c8;
    wire stage0_r48_c7;
    wire stage0_r49_c6;
    wire stage0_r50_c5;
    wire stage0_r51_c4;
    wire stage0_r52_c3;
    wire stage0_r53_c2;
    wire stage0_r54_c1;
    wire stage0_r55_c0;
    wire stage0_r16_c40;
    wire stage0_r17_c39;
    wire stage0_r18_c38;
    wire stage0_r19_c37;
    wire stage0_r20_c36;
    wire stage0_r21_c35;
    wire stage0_r22_c34;
    wire stage0_r23_c33;
    wire stage0_r24_c32;
    wire stage0_r25_c31;
    wire stage0_r26_c30;
    wire stage0_r27_c29;
    wire stage0_r28_c28;
    wire stage0_r29_c27;
    wire stage0_r30_c26;
    wire stage0_r31_c25;
    wire stage0_r32_c24;
    wire stage0_r33_c23;
    wire stage0_r34_c22;
    wire stage0_r35_c21;
    wire stage0_r36_c20;
    wire stage0_r37_c19;
    wire stage0_r38_c18;
    wire stage0_r39_c17;
    wire stage0_r40_c16;
    wire stage0_r41_c15;
    wire stage0_r42_c14;
    wire stage0_r43_c13;
    wire stage0_r44_c12;
    wire stage0_r45_c11;
    wire stage0_r46_c10;
    wire stage0_r47_c9;
    wire stage0_r48_c8;
    wire stage0_r49_c7;
    wire stage0_r50_c6;
    wire stage0_r51_c5;
    wire stage0_r52_c4;
    wire stage0_r53_c3;
    wire stage0_r54_c2;
    wire stage0_r55_c1;
    wire stage0_r56_c0;
    wire stage0_r17_c40;
    wire stage0_r18_c39;
    wire stage0_r19_c38;
    wire stage0_r20_c37;
    wire stage0_r21_c36;
    wire stage0_r22_c35;
    wire stage0_r23_c34;
    wire stage0_r24_c33;
    wire stage0_r25_c32;
    wire stage0_r26_c31;
    wire stage0_r27_c30;
    wire stage0_r28_c29;
    wire stage0_r29_c28;
    wire stage0_r30_c27;
    wire stage0_r31_c26;
    wire stage0_r32_c25;
    wire stage0_r33_c24;
    wire stage0_r34_c23;
    wire stage0_r35_c22;
    wire stage0_r36_c21;
    wire stage0_r37_c20;
    wire stage0_r38_c19;
    wire stage0_r39_c18;
    wire stage0_r40_c17;
    wire stage0_r41_c16;
    wire stage0_r42_c15;
    wire stage0_r43_c14;
    wire stage0_r44_c13;
    wire stage0_r45_c12;
    wire stage0_r46_c11;
    wire stage0_r47_c10;
    wire stage0_r48_c9;
    wire stage0_r49_c8;
    wire stage0_r50_c7;
    wire stage0_r51_c6;
    wire stage0_r52_c5;
    wire stage0_r53_c4;
    wire stage0_r54_c3;
    wire stage0_r55_c2;
    wire stage0_r56_c1;
    wire stage0_r57_c0;
    wire stage0_r18_c40;
    wire stage0_r19_c39;
    wire stage0_r20_c38;
    wire stage0_r21_c37;
    wire stage0_r22_c36;
    wire stage0_r23_c35;
    wire stage0_r24_c34;
    wire stage0_r25_c33;
    wire stage0_r26_c32;
    wire stage0_r27_c31;
    wire stage0_r28_c30;
    wire stage0_r29_c29;
    wire stage0_r30_c28;
    wire stage0_r31_c27;
    wire stage0_r32_c26;
    wire stage0_r33_c25;
    wire stage0_r34_c24;
    wire stage0_r35_c23;
    wire stage0_r36_c22;
    wire stage0_r37_c21;
    wire stage0_r38_c20;
    wire stage0_r39_c19;
    wire stage0_r40_c18;
    wire stage0_r41_c17;
    wire stage0_r42_c16;
    wire stage0_r43_c15;
    wire stage0_r44_c14;
    wire stage0_r45_c13;
    wire stage0_r46_c12;
    wire stage0_r47_c11;
    wire stage0_r48_c10;
    wire stage0_r49_c9;
    wire stage0_r50_c8;
    wire stage0_r51_c7;
    wire stage0_r52_c6;
    wire stage0_r53_c5;
    wire stage0_r54_c4;
    wire stage0_r55_c3;
    wire stage0_r56_c2;
    wire stage0_r57_c1;
    wire stage0_r58_c0;
    wire stage0_r19_c40;
    wire stage0_r20_c39;
    wire stage0_r21_c38;
    wire stage0_r22_c37;
    wire stage0_r23_c36;
    wire stage0_r24_c35;
    wire stage0_r25_c34;
    wire stage0_r26_c33;
    wire stage0_r27_c32;
    wire stage0_r28_c31;
    wire stage0_r29_c30;
    wire stage0_r30_c29;
    wire stage0_r31_c28;
    wire stage0_r32_c27;
    wire stage0_r33_c26;
    wire stage0_r34_c25;
    wire stage0_r35_c24;
    wire stage0_r36_c23;
    wire stage0_r37_c22;
    wire stage0_r38_c21;
    wire stage0_r39_c20;
    wire stage0_r40_c19;
    wire stage0_r41_c18;
    wire stage0_r42_c17;
    wire stage0_r43_c16;
    wire stage0_r44_c15;
    wire stage0_r45_c14;
    wire stage0_r46_c13;
    wire stage0_r47_c12;
    wire stage0_r48_c11;
    wire stage0_r49_c10;
    wire stage0_r50_c9;
    wire stage0_r51_c8;
    wire stage0_r52_c7;
    wire stage0_r53_c6;
    wire stage0_r54_c5;
    wire stage0_r55_c4;
    wire stage0_r56_c3;
    wire stage0_r57_c2;
    wire stage0_r58_c1;
    wire stage0_r59_c0;
    wire stage0_r20_c40;
    wire stage0_r21_c39;
    wire stage0_r22_c38;
    wire stage0_r23_c37;
    wire stage0_r24_c36;
    wire stage0_r25_c35;
    wire stage0_r26_c34;
    wire stage0_r27_c33;
    wire stage0_r28_c32;
    wire stage0_r29_c31;
    wire stage0_r30_c30;
    wire stage0_r31_c29;
    wire stage0_r32_c28;
    wire stage0_r33_c27;
    wire stage0_r34_c26;
    wire stage0_r35_c25;
    wire stage0_r36_c24;
    wire stage0_r37_c23;
    wire stage0_r38_c22;
    wire stage0_r39_c21;
    wire stage0_r40_c20;
    wire stage0_r41_c19;
    wire stage0_r42_c18;
    wire stage0_r43_c17;
    wire stage0_r44_c16;
    wire stage0_r45_c15;
    wire stage0_r46_c14;
    wire stage0_r47_c13;
    wire stage0_r48_c12;
    wire stage0_r49_c11;
    wire stage0_r50_c10;
    wire stage0_r51_c9;
    wire stage0_r52_c8;
    wire stage0_r53_c7;
    wire stage0_r54_c6;
    wire stage0_r55_c5;
    wire stage0_r56_c4;
    wire stage0_r57_c3;
    wire stage0_r58_c2;
    wire stage0_r59_c1;
    wire stage0_r60_c0;
    wire stage0_r21_c40;
    wire stage0_r22_c39;
    wire stage0_r23_c38;
    wire stage0_r24_c37;
    wire stage0_r25_c36;
    wire stage0_r26_c35;
    wire stage0_r27_c34;
    wire stage0_r28_c33;
    wire stage0_r29_c32;
    wire stage0_r30_c31;
    wire stage0_r31_c30;
    wire stage0_r32_c29;
    wire stage0_r33_c28;
    wire stage0_r34_c27;
    wire stage0_r35_c26;
    wire stage0_r36_c25;
    wire stage0_r37_c24;
    wire stage0_r38_c23;
    wire stage0_r39_c22;
    wire stage0_r40_c21;
    wire stage0_r41_c20;
    wire stage0_r42_c19;
    wire stage0_r43_c18;
    wire stage0_r44_c17;
    wire stage0_r45_c16;
    wire stage0_r46_c15;
    wire stage0_r47_c14;
    wire stage0_r48_c13;
    wire stage0_r49_c12;
    wire stage0_r50_c11;
    wire stage0_r51_c10;
    wire stage0_r52_c9;
    wire stage0_r53_c8;
    wire stage0_r54_c7;
    wire stage0_r55_c6;
    wire stage0_r56_c5;
    wire stage0_r57_c4;
    wire stage0_r58_c3;
    wire stage0_r59_c2;
    wire stage0_r60_c1;
    wire stage0_r61_c0;
    wire stage0_r22_c40;
    wire stage0_r23_c39;
    wire stage0_r24_c38;
    wire stage0_r25_c37;
    wire stage0_r26_c36;
    wire stage0_r27_c35;
    wire stage0_r28_c34;
    wire stage0_r29_c33;
    wire stage0_r30_c32;
    wire stage0_r31_c31;
    wire stage0_r32_c30;
    wire stage0_r33_c29;
    wire stage0_r34_c28;
    wire stage0_r35_c27;
    wire stage0_r36_c26;
    wire stage0_r37_c25;
    wire stage0_r38_c24;
    wire stage0_r39_c23;
    wire stage0_r40_c22;
    wire stage0_r41_c21;
    wire stage0_r42_c20;
    wire stage0_r43_c19;
    wire stage0_r44_c18;
    wire stage0_r45_c17;
    wire stage0_r46_c16;
    wire stage0_r47_c15;
    wire stage0_r48_c14;
    wire stage0_r49_c13;
    wire stage0_r50_c12;
    wire stage0_r51_c11;
    wire stage0_r52_c10;
    wire stage0_r53_c9;
    wire stage0_r54_c8;
    wire stage0_r55_c7;
    wire stage0_r56_c6;
    wire stage0_r57_c5;
    wire stage0_r58_c4;
    wire stage0_r59_c3;
    wire stage0_r60_c2;
    wire stage0_r61_c1;
    wire stage0_r62_c0;
    wire stage0_r23_c40;
    wire stage0_r24_c39;
    wire stage0_r25_c38;
    wire stage0_r26_c37;
    wire stage0_r27_c36;
    wire stage0_r28_c35;
    wire stage0_r29_c34;
    wire stage0_r30_c33;
    wire stage0_r31_c32;
    wire stage0_r32_c31;
    wire stage0_r33_c30;
    wire stage0_r34_c29;
    wire stage0_r35_c28;
    wire stage0_r36_c27;
    wire stage0_r37_c26;
    wire stage0_r38_c25;
    wire stage0_r39_c24;
    wire stage0_r40_c23;
    wire stage0_r41_c22;
    wire stage0_r42_c21;
    wire stage0_r43_c20;
    wire stage0_r44_c19;
    wire stage0_r45_c18;
    wire stage0_r46_c17;
    wire stage0_r47_c16;
    wire stage0_r48_c15;
    wire stage0_r49_c14;
    wire stage0_r50_c13;
    wire stage0_r51_c12;
    wire stage0_r52_c11;
    wire stage0_r53_c10;
    wire stage0_r54_c9;
    wire stage0_r55_c8;
    wire stage0_r56_c7;
    wire stage0_r57_c6;
    wire stage0_r58_c5;
    wire stage0_r59_c4;
    wire stage0_r60_c3;
    wire stage0_r61_c2;
    wire stage0_r62_c1;
    wire stage0_r63_c0;
    wire stage0_r24_c40;
    wire stage0_r25_c39;
    wire stage0_r26_c38;
    wire stage0_r27_c37;
    wire stage0_r28_c36;
    wire stage0_r29_c35;
    wire stage0_r30_c34;
    wire stage0_r31_c33;
    wire stage0_r32_c32;
    wire stage0_r33_c31;
    wire stage0_r34_c30;
    wire stage0_r35_c29;
    wire stage0_r36_c28;
    wire stage0_r37_c27;
    wire stage0_r38_c26;
    wire stage0_r39_c25;
    wire stage0_r40_c24;
    wire stage0_r41_c23;
    wire stage0_r42_c22;
    wire stage0_r43_c21;
    wire stage0_r44_c20;
    wire stage0_r45_c19;
    wire stage0_r46_c18;
    wire stage0_r47_c17;
    wire stage0_r48_c16;
    wire stage0_r49_c15;
    wire stage0_r50_c14;
    wire stage0_r51_c13;
    wire stage0_r52_c12;
    wire stage0_r53_c11;
    wire stage0_r54_c10;
    wire stage0_r55_c9;
    wire stage0_r56_c8;
    wire stage0_r57_c7;
    wire stage0_r58_c6;
    wire stage0_r59_c5;
    wire stage0_r60_c4;
    wire stage0_r61_c3;
    wire stage0_r62_c2;
    wire stage0_r63_c1;
    wire stage0_r64_c0;
    wire stage0_r25_c40;
    wire stage0_r26_c39;
    wire stage0_r27_c38;
    wire stage0_r28_c37;
    wire stage0_r29_c36;
    wire stage0_r30_c35;
    wire stage0_r31_c34;
    wire stage0_r32_c33;
    wire stage0_r33_c32;
    wire stage0_r34_c31;
    wire stage0_r35_c30;
    wire stage0_r36_c29;
    wire stage0_r37_c28;
    wire stage0_r38_c27;
    wire stage0_r39_c26;
    wire stage0_r40_c25;
    wire stage0_r41_c24;
    wire stage0_r42_c23;
    wire stage0_r43_c22;
    wire stage0_r44_c21;
    wire stage0_r45_c20;
    wire stage0_r46_c19;
    wire stage0_r47_c18;
    wire stage0_r48_c17;
    wire stage0_r49_c16;
    wire stage0_r50_c15;
    wire stage0_r51_c14;
    wire stage0_r52_c13;
    wire stage0_r53_c12;
    wire stage0_r54_c11;
    wire stage0_r55_c10;
    wire stage0_r56_c9;
    wire stage0_r57_c8;
    wire stage0_r58_c7;
    wire stage0_r59_c6;
    wire stage0_r60_c5;
    wire stage0_r61_c4;
    wire stage0_r62_c3;
    wire stage0_r63_c2;
    wire stage0_r64_c1;
    wire stage0_r65_c0;
    wire stage0_r26_c40;
    wire stage0_r27_c39;
    wire stage0_r28_c38;
    wire stage0_r29_c37;
    wire stage0_r30_c36;
    wire stage0_r31_c35;
    wire stage0_r32_c34;
    wire stage0_r33_c33;
    wire stage0_r34_c32;
    wire stage0_r35_c31;
    wire stage0_r36_c30;
    wire stage0_r37_c29;
    wire stage0_r38_c28;
    wire stage0_r39_c27;
    wire stage0_r40_c26;
    wire stage0_r41_c25;
    wire stage0_r42_c24;
    wire stage0_r43_c23;
    wire stage0_r44_c22;
    wire stage0_r45_c21;
    wire stage0_r46_c20;
    wire stage0_r47_c19;
    wire stage0_r48_c18;
    wire stage0_r49_c17;
    wire stage0_r50_c16;
    wire stage0_r51_c15;
    wire stage0_r52_c14;
    wire stage0_r53_c13;
    wire stage0_r54_c12;
    wire stage0_r55_c11;
    wire stage0_r56_c10;
    wire stage0_r57_c9;
    wire stage0_r58_c8;
    wire stage0_r59_c7;
    wire stage0_r60_c6;
    wire stage0_r61_c5;
    wire stage0_r62_c4;
    wire stage0_r63_c3;
    wire stage0_r64_c2;
    wire stage0_r65_c1;
    wire stage0_r66_c0;
    wire stage0_r27_c40;
    wire stage0_r28_c39;
    wire stage0_r29_c38;
    wire stage0_r30_c37;
    wire stage0_r31_c36;
    wire stage0_r32_c35;
    wire stage0_r33_c34;
    wire stage0_r34_c33;
    wire stage0_r35_c32;
    wire stage0_r36_c31;
    wire stage0_r37_c30;
    wire stage0_r38_c29;
    wire stage0_r39_c28;
    wire stage0_r40_c27;
    wire stage0_r41_c26;
    wire stage0_r42_c25;
    wire stage0_r43_c24;
    wire stage0_r44_c23;
    wire stage0_r45_c22;
    wire stage0_r46_c21;
    wire stage0_r47_c20;
    wire stage0_r48_c19;
    wire stage0_r49_c18;
    wire stage0_r50_c17;
    wire stage0_r51_c16;
    wire stage0_r52_c15;
    wire stage0_r53_c14;
    wire stage0_r54_c13;
    wire stage0_r55_c12;
    wire stage0_r56_c11;
    wire stage0_r57_c10;
    wire stage0_r58_c9;
    wire stage0_r59_c8;
    wire stage0_r60_c7;
    wire stage0_r61_c6;
    wire stage0_r62_c5;
    wire stage0_r63_c4;
    wire stage0_r64_c3;
    wire stage0_r65_c2;
    wire stage0_r66_c1;
    wire stage0_r67_c0;
    wire stage0_r28_c40;
    wire stage0_r29_c39;
    wire stage0_r30_c38;
    wire stage0_r31_c37;
    wire stage0_r32_c36;
    wire stage0_r33_c35;
    wire stage0_r34_c34;
    wire stage0_r35_c33;
    wire stage0_r36_c32;
    wire stage0_r37_c31;
    wire stage0_r38_c30;
    wire stage0_r39_c29;
    wire stage0_r40_c28;
    wire stage0_r41_c27;
    wire stage0_r42_c26;
    wire stage0_r43_c25;
    wire stage0_r44_c24;
    wire stage0_r45_c23;
    wire stage0_r46_c22;
    wire stage0_r47_c21;
    wire stage0_r48_c20;
    wire stage0_r49_c19;
    wire stage0_r50_c18;
    wire stage0_r51_c17;
    wire stage0_r52_c16;
    wire stage0_r53_c15;
    wire stage0_r54_c14;
    wire stage0_r55_c13;
    wire stage0_r56_c12;
    wire stage0_r57_c11;
    wire stage0_r58_c10;
    wire stage0_r59_c9;
    wire stage0_r60_c8;
    wire stage0_r61_c7;
    wire stage0_r62_c6;
    wire stage0_r63_c5;
    wire stage0_r64_c4;
    wire stage0_r65_c3;
    wire stage0_r66_c2;
    wire stage0_r67_c1;
    wire stage0_r68_c0;
    wire stage0_r29_c40;
    wire stage0_r30_c39;
    wire stage0_r31_c38;
    wire stage0_r32_c37;
    wire stage0_r33_c36;
    wire stage0_r34_c35;
    wire stage0_r35_c34;
    wire stage0_r36_c33;
    wire stage0_r37_c32;
    wire stage0_r38_c31;
    wire stage0_r39_c30;
    wire stage0_r40_c29;
    wire stage0_r41_c28;
    wire stage0_r42_c27;
    wire stage0_r43_c26;
    wire stage0_r44_c25;
    wire stage0_r45_c24;
    wire stage0_r46_c23;
    wire stage0_r47_c22;
    wire stage0_r48_c21;
    wire stage0_r49_c20;
    wire stage0_r50_c19;
    wire stage0_r51_c18;
    wire stage0_r52_c17;
    wire stage0_r53_c16;
    wire stage0_r54_c15;
    wire stage0_r55_c14;
    wire stage0_r56_c13;
    wire stage0_r57_c12;
    wire stage0_r58_c11;
    wire stage0_r59_c10;
    wire stage0_r60_c9;
    wire stage0_r61_c8;
    wire stage0_r62_c7;
    wire stage0_r63_c6;
    wire stage0_r64_c5;
    wire stage0_r65_c4;
    wire stage0_r66_c3;
    wire stage0_r67_c2;
    wire stage0_r68_c1;
    wire stage0_r69_c0;
    wire stage0_r30_c40;
    wire stage0_r31_c39;
    wire stage0_r32_c38;
    wire stage0_r33_c37;
    wire stage0_r34_c36;
    wire stage0_r35_c35;
    wire stage0_r36_c34;
    wire stage0_r37_c33;
    wire stage0_r38_c32;
    wire stage0_r39_c31;
    wire stage0_r40_c30;
    wire stage0_r41_c29;
    wire stage0_r42_c28;
    wire stage0_r43_c27;
    wire stage0_r44_c26;
    wire stage0_r45_c25;
    wire stage0_r46_c24;
    wire stage0_r47_c23;
    wire stage0_r48_c22;
    wire stage0_r49_c21;
    wire stage0_r50_c20;
    wire stage0_r51_c19;
    wire stage0_r52_c18;
    wire stage0_r53_c17;
    wire stage0_r54_c16;
    wire stage0_r55_c15;
    wire stage0_r56_c14;
    wire stage0_r57_c13;
    wire stage0_r58_c12;
    wire stage0_r59_c11;
    wire stage0_r60_c10;
    wire stage0_r61_c9;
    wire stage0_r62_c8;
    wire stage0_r63_c7;
    wire stage0_r64_c6;
    wire stage0_r65_c5;
    wire stage0_r66_c4;
    wire stage0_r67_c3;
    wire stage0_r68_c2;
    wire stage0_r69_c1;
    wire stage0_r70_c0;
    wire stage0_r31_c40;
    wire stage0_r32_c39;
    wire stage0_r33_c38;
    wire stage0_r34_c37;
    wire stage0_r35_c36;
    wire stage0_r36_c35;
    wire stage0_r37_c34;
    wire stage0_r38_c33;
    wire stage0_r39_c32;
    wire stage0_r40_c31;
    wire stage0_r41_c30;
    wire stage0_r42_c29;
    wire stage0_r43_c28;
    wire stage0_r44_c27;
    wire stage0_r45_c26;
    wire stage0_r46_c25;
    wire stage0_r47_c24;
    wire stage0_r48_c23;
    wire stage0_r49_c22;
    wire stage0_r50_c21;
    wire stage0_r51_c20;
    wire stage0_r52_c19;
    wire stage0_r53_c18;
    wire stage0_r54_c17;
    wire stage0_r55_c16;
    wire stage0_r56_c15;
    wire stage0_r57_c14;
    wire stage0_r58_c13;
    wire stage0_r59_c12;
    wire stage0_r60_c11;
    wire stage0_r61_c10;
    wire stage0_r62_c9;
    wire stage0_r63_c8;
    wire stage0_r64_c7;
    wire stage0_r65_c6;
    wire stage0_r66_c5;
    wire stage0_r67_c4;
    wire stage0_r68_c3;
    wire stage0_r69_c2;
    wire stage0_r70_c1;
    wire stage0_r71_c0;
    wire stage0_r32_c40;
    wire stage0_r33_c39;
    wire stage0_r34_c38;
    wire stage0_r35_c37;
    wire stage0_r36_c36;
    wire stage0_r37_c35;
    wire stage0_r38_c34;
    wire stage0_r39_c33;
    wire stage0_r40_c32;
    wire stage0_r41_c31;
    wire stage0_r42_c30;
    wire stage0_r43_c29;
    wire stage0_r44_c28;
    wire stage0_r45_c27;
    wire stage0_r46_c26;
    wire stage0_r47_c25;
    wire stage0_r48_c24;
    wire stage0_r49_c23;
    wire stage0_r50_c22;
    wire stage0_r51_c21;
    wire stage0_r52_c20;
    wire stage0_r53_c19;
    wire stage0_r54_c18;
    wire stage0_r55_c17;
    wire stage0_r56_c16;
    wire stage0_r57_c15;
    wire stage0_r58_c14;
    wire stage0_r59_c13;
    wire stage0_r60_c12;
    wire stage0_r61_c11;
    wire stage0_r62_c10;
    wire stage0_r63_c9;
    wire stage0_r64_c8;
    wire stage0_r65_c7;
    wire stage0_r66_c6;
    wire stage0_r67_c5;
    wire stage0_r68_c4;
    wire stage0_r69_c3;
    wire stage0_r70_c2;
    wire stage0_r71_c1;
    wire stage0_r33_c40;
    wire stage0_r34_c39;
    wire stage0_r35_c38;
    wire stage0_r36_c37;
    wire stage0_r37_c36;
    wire stage0_r38_c35;
    wire stage0_r39_c34;
    wire stage0_r40_c33;
    wire stage0_r41_c32;
    wire stage0_r42_c31;
    wire stage0_r43_c30;
    wire stage0_r44_c29;
    wire stage0_r45_c28;
    wire stage0_r46_c27;
    wire stage0_r47_c26;
    wire stage0_r48_c25;
    wire stage0_r49_c24;
    wire stage0_r50_c23;
    wire stage0_r51_c22;
    wire stage0_r52_c21;
    wire stage0_r53_c20;
    wire stage0_r54_c19;
    wire stage0_r55_c18;
    wire stage0_r56_c17;
    wire stage0_r57_c16;
    wire stage0_r58_c15;
    wire stage0_r59_c14;
    wire stage0_r60_c13;
    wire stage0_r61_c12;
    wire stage0_r62_c11;
    wire stage0_r63_c10;
    wire stage0_r64_c9;
    wire stage0_r65_c8;
    wire stage0_r66_c7;
    wire stage0_r67_c6;
    wire stage0_r68_c5;
    wire stage0_r69_c4;
    wire stage0_r70_c3;
    wire stage0_r71_c2;
    wire stage0_r34_c40;
    wire stage0_r35_c39;
    wire stage0_r36_c38;
    wire stage0_r37_c37;
    wire stage0_r38_c36;
    wire stage0_r39_c35;
    wire stage0_r40_c34;
    wire stage0_r41_c33;
    wire stage0_r42_c32;
    wire stage0_r43_c31;
    wire stage0_r44_c30;
    wire stage0_r45_c29;
    wire stage0_r46_c28;
    wire stage0_r47_c27;
    wire stage0_r48_c26;
    wire stage0_r49_c25;
    wire stage0_r50_c24;
    wire stage0_r51_c23;
    wire stage0_r52_c22;
    wire stage0_r53_c21;
    wire stage0_r54_c20;
    wire stage0_r55_c19;
    wire stage0_r56_c18;
    wire stage0_r57_c17;
    wire stage0_r58_c16;
    wire stage0_r59_c15;
    wire stage0_r60_c14;
    wire stage0_r61_c13;
    wire stage0_r62_c12;
    wire stage0_r63_c11;
    wire stage0_r64_c10;
    wire stage0_r65_c9;
    wire stage0_r66_c8;
    wire stage0_r67_c7;
    wire stage0_r68_c6;
    wire stage0_r69_c5;
    wire stage0_r70_c4;
    wire stage0_r71_c3;
    wire stage0_r35_c40;
    wire stage0_r36_c39;
    wire stage0_r37_c38;
    wire stage0_r38_c37;
    wire stage0_r39_c36;
    wire stage0_r40_c35;
    wire stage0_r41_c34;
    wire stage0_r42_c33;
    wire stage0_r43_c32;
    wire stage0_r44_c31;
    wire stage0_r45_c30;
    wire stage0_r46_c29;
    wire stage0_r47_c28;
    wire stage0_r48_c27;
    wire stage0_r49_c26;
    wire stage0_r50_c25;
    wire stage0_r51_c24;
    wire stage0_r52_c23;
    wire stage0_r53_c22;
    wire stage0_r54_c21;
    wire stage0_r55_c20;
    wire stage0_r56_c19;
    wire stage0_r57_c18;
    wire stage0_r58_c17;
    wire stage0_r59_c16;
    wire stage0_r60_c15;
    wire stage0_r61_c14;
    wire stage0_r62_c13;
    wire stage0_r63_c12;
    wire stage0_r64_c11;
    wire stage0_r65_c10;
    wire stage0_r66_c9;
    wire stage0_r67_c8;
    wire stage0_r68_c7;
    wire stage0_r69_c6;
    wire stage0_r70_c5;
    wire stage0_r71_c4;
    wire stage0_r36_c40;
    wire stage0_r37_c39;
    wire stage0_r38_c38;
    wire stage0_r39_c37;
    wire stage0_r40_c36;
    wire stage0_r41_c35;
    wire stage0_r42_c34;
    wire stage0_r43_c33;
    wire stage0_r44_c32;
    wire stage0_r45_c31;
    wire stage0_r46_c30;
    wire stage0_r47_c29;
    wire stage0_r48_c28;
    wire stage0_r49_c27;
    wire stage0_r50_c26;
    wire stage0_r51_c25;
    wire stage0_r52_c24;
    wire stage0_r53_c23;
    wire stage0_r54_c22;
    wire stage0_r55_c21;
    wire stage0_r56_c20;
    wire stage0_r57_c19;
    wire stage0_r58_c18;
    wire stage0_r59_c17;
    wire stage0_r60_c16;
    wire stage0_r61_c15;
    wire stage0_r62_c14;
    wire stage0_r63_c13;
    wire stage0_r64_c12;
    wire stage0_r65_c11;
    wire stage0_r66_c10;
    wire stage0_r67_c9;
    wire stage0_r68_c8;
    wire stage0_r69_c7;
    wire stage0_r70_c6;
    wire stage0_r71_c5;
    wire stage0_r37_c40;
    wire stage0_r38_c39;
    wire stage0_r39_c38;
    wire stage0_r40_c37;
    wire stage0_r41_c36;
    wire stage0_r42_c35;
    wire stage0_r43_c34;
    wire stage0_r44_c33;
    wire stage0_r45_c32;
    wire stage0_r46_c31;
    wire stage0_r47_c30;
    wire stage0_r48_c29;
    wire stage0_r49_c28;
    wire stage0_r50_c27;
    wire stage0_r51_c26;
    wire stage0_r52_c25;
    wire stage0_r53_c24;
    wire stage0_r54_c23;
    wire stage0_r55_c22;
    wire stage0_r56_c21;
    wire stage0_r57_c20;
    wire stage0_r58_c19;
    wire stage0_r59_c18;
    wire stage0_r60_c17;
    wire stage0_r61_c16;
    wire stage0_r62_c15;
    wire stage0_r63_c14;
    wire stage0_r64_c13;
    wire stage0_r65_c12;
    wire stage0_r66_c11;
    wire stage0_r67_c10;
    wire stage0_r68_c9;
    wire stage0_r69_c8;
    wire stage0_r70_c7;
    wire stage0_r71_c6;
    wire stage0_r38_c40;
    wire stage0_r39_c39;
    wire stage0_r40_c38;
    wire stage0_r41_c37;
    wire stage0_r42_c36;
    wire stage0_r43_c35;
    wire stage0_r44_c34;
    wire stage0_r45_c33;
    wire stage0_r46_c32;
    wire stage0_r47_c31;
    wire stage0_r48_c30;
    wire stage0_r49_c29;
    wire stage0_r50_c28;
    wire stage0_r51_c27;
    wire stage0_r52_c26;
    wire stage0_r53_c25;
    wire stage0_r54_c24;
    wire stage0_r55_c23;
    wire stage0_r56_c22;
    wire stage0_r57_c21;
    wire stage0_r58_c20;
    wire stage0_r59_c19;
    wire stage0_r60_c18;
    wire stage0_r61_c17;
    wire stage0_r62_c16;
    wire stage0_r63_c15;
    wire stage0_r64_c14;
    wire stage0_r65_c13;
    wire stage0_r66_c12;
    wire stage0_r67_c11;
    wire stage0_r68_c10;
    wire stage0_r69_c9;
    wire stage0_r70_c8;
    wire stage0_r71_c7;
    wire stage0_r39_c40;
    wire stage0_r40_c39;
    wire stage0_r41_c38;
    wire stage0_r42_c37;
    wire stage0_r43_c36;
    wire stage0_r44_c35;
    wire stage0_r45_c34;
    wire stage0_r46_c33;
    wire stage0_r47_c32;
    wire stage0_r48_c31;
    wire stage0_r49_c30;
    wire stage0_r50_c29;
    wire stage0_r51_c28;
    wire stage0_r52_c27;
    wire stage0_r53_c26;
    wire stage0_r54_c25;
    wire stage0_r55_c24;
    wire stage0_r56_c23;
    wire stage0_r57_c22;
    wire stage0_r58_c21;
    wire stage0_r59_c20;
    wire stage0_r60_c19;
    wire stage0_r61_c18;
    wire stage0_r62_c17;
    wire stage0_r63_c16;
    wire stage0_r64_c15;
    wire stage0_r65_c14;
    wire stage0_r66_c13;
    wire stage0_r67_c12;
    wire stage0_r68_c11;
    wire stage0_r69_c10;
    wire stage0_r70_c9;
    wire stage0_r71_c8;
    wire stage0_r40_c40;
    wire stage0_r41_c39;
    wire stage0_r42_c38;
    wire stage0_r43_c37;
    wire stage0_r44_c36;
    wire stage0_r45_c35;
    wire stage0_r46_c34;
    wire stage0_r47_c33;
    wire stage0_r48_c32;
    wire stage0_r49_c31;
    wire stage0_r50_c30;
    wire stage0_r51_c29;
    wire stage0_r52_c28;
    wire stage0_r53_c27;
    wire stage0_r54_c26;
    wire stage0_r55_c25;
    wire stage0_r56_c24;
    wire stage0_r57_c23;
    wire stage0_r58_c22;
    wire stage0_r59_c21;
    wire stage0_r60_c20;
    wire stage0_r61_c19;
    wire stage0_r62_c18;
    wire stage0_r63_c17;
    wire stage0_r64_c16;
    wire stage0_r65_c15;
    wire stage0_r66_c14;
    wire stage0_r67_c13;
    wire stage0_r68_c12;
    wire stage0_r69_c11;
    wire stage0_r70_c10;
    wire stage0_r71_c9;
    wire stage0_r41_c40;
    wire stage0_r42_c39;
    wire stage0_r43_c38;
    wire stage0_r44_c37;
    wire stage0_r45_c36;
    wire stage0_r46_c35;
    wire stage0_r47_c34;
    wire stage0_r48_c33;
    wire stage0_r49_c32;
    wire stage0_r50_c31;
    wire stage0_r51_c30;
    wire stage0_r52_c29;
    wire stage0_r53_c28;
    wire stage0_r54_c27;
    wire stage0_r55_c26;
    wire stage0_r56_c25;
    wire stage0_r57_c24;
    wire stage0_r58_c23;
    wire stage0_r59_c22;
    wire stage0_r60_c21;
    wire stage0_r61_c20;
    wire stage0_r62_c19;
    wire stage0_r63_c18;
    wire stage0_r64_c17;
    wire stage0_r65_c16;
    wire stage0_r66_c15;
    wire stage0_r67_c14;
    wire stage0_r68_c13;
    wire stage0_r69_c12;
    wire stage0_r70_c11;
    wire stage0_r71_c10;
    wire stage0_r42_c40;
    wire stage0_r43_c39;
    wire stage0_r44_c38;
    wire stage0_r45_c37;
    wire stage0_r46_c36;
    wire stage0_r47_c35;
    wire stage0_r48_c34;
    wire stage0_r49_c33;
    wire stage0_r50_c32;
    wire stage0_r51_c31;
    wire stage0_r52_c30;
    wire stage0_r53_c29;
    wire stage0_r54_c28;
    wire stage0_r55_c27;
    wire stage0_r56_c26;
    wire stage0_r57_c25;
    wire stage0_r58_c24;
    wire stage0_r59_c23;
    wire stage0_r60_c22;
    wire stage0_r61_c21;
    wire stage0_r62_c20;
    wire stage0_r63_c19;
    wire stage0_r64_c18;
    wire stage0_r65_c17;
    wire stage0_r66_c16;
    wire stage0_r67_c15;
    wire stage0_r68_c14;
    wire stage0_r69_c13;
    wire stage0_r70_c12;
    wire stage0_r71_c11;
    wire stage0_r43_c40;
    wire stage0_r44_c39;
    wire stage0_r45_c38;
    wire stage0_r46_c37;
    wire stage0_r47_c36;
    wire stage0_r48_c35;
    wire stage0_r49_c34;
    wire stage0_r50_c33;
    wire stage0_r51_c32;
    wire stage0_r52_c31;
    wire stage0_r53_c30;
    wire stage0_r54_c29;
    wire stage0_r55_c28;
    wire stage0_r56_c27;
    wire stage0_r57_c26;
    wire stage0_r58_c25;
    wire stage0_r59_c24;
    wire stage0_r60_c23;
    wire stage0_r61_c22;
    wire stage0_r62_c21;
    wire stage0_r63_c20;
    wire stage0_r64_c19;
    wire stage0_r65_c18;
    wire stage0_r66_c17;
    wire stage0_r67_c16;
    wire stage0_r68_c15;
    wire stage0_r69_c14;
    wire stage0_r70_c13;
    wire stage0_r71_c12;
    wire stage0_r44_c40;
    wire stage0_r45_c39;
    wire stage0_r46_c38;
    wire stage0_r47_c37;
    wire stage0_r48_c36;
    wire stage0_r49_c35;
    wire stage0_r50_c34;
    wire stage0_r51_c33;
    wire stage0_r52_c32;
    wire stage0_r53_c31;
    wire stage0_r54_c30;
    wire stage0_r55_c29;
    wire stage0_r56_c28;
    wire stage0_r57_c27;
    wire stage0_r58_c26;
    wire stage0_r59_c25;
    wire stage0_r60_c24;
    wire stage0_r61_c23;
    wire stage0_r62_c22;
    wire stage0_r63_c21;
    wire stage0_r64_c20;
    wire stage0_r65_c19;
    wire stage0_r66_c18;
    wire stage0_r67_c17;
    wire stage0_r68_c16;
    wire stage0_r69_c15;
    wire stage0_r70_c14;
    wire stage0_r71_c13;
    wire stage0_r45_c40;
    wire stage0_r46_c39;
    wire stage0_r47_c38;
    wire stage0_r48_c37;
    wire stage0_r49_c36;
    wire stage0_r50_c35;
    wire stage0_r51_c34;
    wire stage0_r52_c33;
    wire stage0_r53_c32;
    wire stage0_r54_c31;
    wire stage0_r55_c30;
    wire stage0_r56_c29;
    wire stage0_r57_c28;
    wire stage0_r58_c27;
    wire stage0_r59_c26;
    wire stage0_r60_c25;
    wire stage0_r61_c24;
    wire stage0_r62_c23;
    wire stage0_r63_c22;
    wire stage0_r64_c21;
    wire stage0_r65_c20;
    wire stage0_r66_c19;
    wire stage0_r67_c18;
    wire stage0_r68_c17;
    wire stage0_r69_c16;
    wire stage0_r70_c15;
    wire stage0_r71_c14;
    wire stage0_r46_c40;
    wire stage0_r47_c39;
    wire stage0_r48_c38;
    wire stage0_r49_c37;
    wire stage0_r50_c36;
    wire stage0_r51_c35;
    wire stage0_r52_c34;
    wire stage0_r53_c33;
    wire stage0_r54_c32;
    wire stage0_r55_c31;
    wire stage0_r56_c30;
    wire stage0_r57_c29;
    wire stage0_r58_c28;
    wire stage0_r59_c27;
    wire stage0_r60_c26;
    wire stage0_r61_c25;
    wire stage0_r62_c24;
    wire stage0_r63_c23;
    wire stage0_r64_c22;
    wire stage0_r65_c21;
    wire stage0_r66_c20;
    wire stage0_r67_c19;
    wire stage0_r68_c18;
    wire stage0_r69_c17;
    wire stage0_r70_c16;
    wire stage0_r71_c15;
    wire stage0_r47_c40;
    wire stage0_r48_c39;
    wire stage0_r49_c38;
    wire stage0_r50_c37;
    wire stage0_r51_c36;
    wire stage0_r52_c35;
    wire stage0_r53_c34;
    wire stage0_r54_c33;
    wire stage0_r55_c32;
    wire stage0_r56_c31;
    wire stage0_r57_c30;
    wire stage0_r58_c29;
    wire stage0_r59_c28;
    wire stage0_r60_c27;
    wire stage0_r61_c26;
    wire stage0_r62_c25;
    wire stage0_r63_c24;
    wire stage0_r64_c23;
    wire stage0_r65_c22;
    wire stage0_r66_c21;
    wire stage0_r67_c20;
    wire stage0_r68_c19;
    wire stage0_r69_c18;
    wire stage0_r70_c17;
    wire stage0_r71_c16;
    wire stage0_r48_c40;
    wire stage0_r49_c39;
    wire stage0_r50_c38;
    wire stage0_r51_c37;
    wire stage0_r52_c36;
    wire stage0_r53_c35;
    wire stage0_r54_c34;
    wire stage0_r55_c33;
    wire stage0_r56_c32;
    wire stage0_r57_c31;
    wire stage0_r58_c30;
    wire stage0_r59_c29;
    wire stage0_r60_c28;
    wire stage0_r61_c27;
    wire stage0_r62_c26;
    wire stage0_r63_c25;
    wire stage0_r64_c24;
    wire stage0_r65_c23;
    wire stage0_r66_c22;
    wire stage0_r67_c21;
    wire stage0_r68_c20;
    wire stage0_r69_c19;
    wire stage0_r70_c18;
    wire stage0_r71_c17;
    wire stage0_r49_c40;
    wire stage0_r50_c39;
    wire stage0_r51_c38;
    wire stage0_r52_c37;
    wire stage0_r53_c36;
    wire stage0_r54_c35;
    wire stage0_r55_c34;
    wire stage0_r56_c33;
    wire stage0_r57_c32;
    wire stage0_r58_c31;
    wire stage0_r59_c30;
    wire stage0_r60_c29;
    wire stage0_r61_c28;
    wire stage0_r62_c27;
    wire stage0_r63_c26;
    wire stage0_r64_c25;
    wire stage0_r65_c24;
    wire stage0_r66_c23;
    wire stage0_r67_c22;
    wire stage0_r68_c21;
    wire stage0_r69_c20;
    wire stage0_r70_c19;
    wire stage0_r71_c18;
    wire stage0_r50_c40;
    wire stage0_r51_c39;
    wire stage0_r52_c38;
    wire stage0_r53_c37;
    wire stage0_r54_c36;
    wire stage0_r55_c35;
    wire stage0_r56_c34;
    wire stage0_r57_c33;
    wire stage0_r58_c32;
    wire stage0_r59_c31;
    wire stage0_r60_c30;
    wire stage0_r61_c29;
    wire stage0_r62_c28;
    wire stage0_r63_c27;
    wire stage0_r64_c26;
    wire stage0_r65_c25;
    wire stage0_r66_c24;
    wire stage0_r67_c23;
    wire stage0_r68_c22;
    wire stage0_r69_c21;
    wire stage0_r70_c20;
    wire stage0_r71_c19;
    wire stage0_r51_c40;
    wire stage0_r52_c39;
    wire stage0_r53_c38;
    wire stage0_r54_c37;
    wire stage0_r55_c36;
    wire stage0_r56_c35;
    wire stage0_r57_c34;
    wire stage0_r58_c33;
    wire stage0_r59_c32;
    wire stage0_r60_c31;
    wire stage0_r61_c30;
    wire stage0_r62_c29;
    wire stage0_r63_c28;
    wire stage0_r64_c27;
    wire stage0_r65_c26;
    wire stage0_r66_c25;
    wire stage0_r67_c24;
    wire stage0_r68_c23;
    wire stage0_r69_c22;
    wire stage0_r70_c21;
    wire stage0_r71_c20;
    wire stage0_r52_c40;
    wire stage0_r53_c39;
    wire stage0_r54_c38;
    wire stage0_r55_c37;
    wire stage0_r56_c36;
    wire stage0_r57_c35;
    wire stage0_r58_c34;
    wire stage0_r59_c33;
    wire stage0_r60_c32;
    wire stage0_r61_c31;
    wire stage0_r62_c30;
    wire stage0_r63_c29;
    wire stage0_r64_c28;
    wire stage0_r65_c27;
    wire stage0_r66_c26;
    wire stage0_r67_c25;
    wire stage0_r68_c24;
    wire stage0_r69_c23;
    wire stage0_r70_c22;
    wire stage0_r71_c21;
    wire stage0_r53_c40;
    wire stage0_r54_c39;
    wire stage0_r55_c38;
    wire stage0_r56_c37;
    wire stage0_r57_c36;
    wire stage0_r58_c35;
    wire stage0_r59_c34;
    wire stage0_r60_c33;
    wire stage0_r61_c32;
    wire stage0_r62_c31;
    wire stage0_r63_c30;
    wire stage0_r64_c29;
    wire stage0_r65_c28;
    wire stage0_r66_c27;
    wire stage0_r67_c26;
    wire stage0_r68_c25;
    wire stage0_r69_c24;
    wire stage0_r70_c23;
    wire stage0_r71_c22;
    wire stage0_r54_c40;
    wire stage0_r55_c39;
    wire stage0_r56_c38;
    wire stage0_r57_c37;
    wire stage0_r58_c36;
    wire stage0_r59_c35;
    wire stage0_r60_c34;
    wire stage0_r61_c33;
    wire stage0_r62_c32;
    wire stage0_r63_c31;
    wire stage0_r64_c30;
    wire stage0_r65_c29;
    wire stage0_r66_c28;
    wire stage0_r67_c27;
    wire stage0_r68_c26;
    wire stage0_r69_c25;
    wire stage0_r70_c24;
    wire stage0_r71_c23;
    wire stage0_r55_c40;
    wire stage0_r56_c39;
    wire stage0_r57_c38;
    wire stage0_r58_c37;
    wire stage0_r59_c36;
    wire stage0_r60_c35;
    wire stage0_r61_c34;
    wire stage0_r62_c33;
    wire stage0_r63_c32;
    wire stage0_r64_c31;
    wire stage0_r65_c30;
    wire stage0_r66_c29;
    wire stage0_r67_c28;
    wire stage0_r68_c27;
    wire stage0_r69_c26;
    wire stage0_r70_c25;
    wire stage0_r71_c24;
    wire stage0_r56_c40;
    wire stage0_r57_c39;
    wire stage0_r58_c38;
    wire stage0_r59_c37;
    wire stage0_r60_c36;
    wire stage0_r61_c35;
    wire stage0_r62_c34;
    wire stage0_r63_c33;
    wire stage0_r64_c32;
    wire stage0_r65_c31;
    wire stage0_r66_c30;
    wire stage0_r67_c29;
    wire stage0_r68_c28;
    wire stage0_r69_c27;
    wire stage0_r70_c26;
    wire stage0_r71_c25;
    wire stage0_r57_c40;
    wire stage0_r58_c39;
    wire stage0_r59_c38;
    wire stage0_r60_c37;
    wire stage0_r61_c36;
    wire stage0_r62_c35;
    wire stage0_r63_c34;
    wire stage0_r64_c33;
    wire stage0_r65_c32;
    wire stage0_r66_c31;
    wire stage0_r67_c30;
    wire stage0_r68_c29;
    wire stage0_r69_c28;
    wire stage0_r70_c27;
    wire stage0_r71_c26;
    wire stage0_r58_c40;
    wire stage0_r59_c39;
    wire stage0_r60_c38;
    wire stage0_r61_c37;
    wire stage0_r62_c36;
    wire stage0_r63_c35;
    wire stage0_r64_c34;
    wire stage0_r65_c33;
    wire stage0_r66_c32;
    wire stage0_r67_c31;
    wire stage0_r68_c30;
    wire stage0_r69_c29;
    wire stage0_r70_c28;
    wire stage0_r71_c27;
    wire stage0_r59_c40;
    wire stage0_r60_c39;
    wire stage0_r61_c38;
    wire stage0_r62_c37;
    wire stage0_r63_c36;
    wire stage0_r64_c35;
    wire stage0_r65_c34;
    wire stage0_r66_c33;
    wire stage0_r67_c32;
    wire stage0_r68_c31;
    wire stage0_r69_c30;
    wire stage0_r70_c29;
    wire stage0_r71_c28;
    wire stage0_r60_c40;
    wire stage0_r61_c39;
    wire stage0_r62_c38;
    wire stage0_r63_c37;
    wire stage0_r64_c36;
    wire stage0_r65_c35;
    wire stage0_r66_c34;
    wire stage0_r67_c33;
    wire stage0_r68_c32;
    wire stage0_r69_c31;
    wire stage0_r70_c30;
    wire stage0_r71_c29;
    wire stage0_r61_c40;
    wire stage0_r62_c39;
    wire stage0_r63_c38;
    wire stage0_r64_c37;
    wire stage0_r65_c36;
    wire stage0_r66_c35;
    wire stage0_r67_c34;
    wire stage0_r68_c33;
    wire stage0_r69_c32;
    wire stage0_r70_c31;
    wire stage0_r71_c30;
    wire stage0_r62_c40;
    wire stage0_r63_c39;
    wire stage0_r64_c38;
    wire stage0_r65_c37;
    wire stage0_r66_c36;
    wire stage0_r67_c35;
    wire stage0_r68_c34;
    wire stage0_r69_c33;
    wire stage0_r70_c32;
    wire stage0_r71_c31;
    wire stage0_r63_c40;
    wire stage0_r64_c39;
    wire stage0_r65_c38;
    wire stage0_r66_c37;
    wire stage0_r67_c36;
    wire stage0_r68_c35;
    wire stage0_r69_c34;
    wire stage0_r70_c33;
    wire stage0_r71_c32;
    wire stage0_r64_c40;
    wire stage0_r65_c39;
    wire stage0_r66_c38;
    wire stage0_r67_c37;
    wire stage0_r68_c36;
    wire stage0_r69_c35;
    wire stage0_r70_c34;
    wire stage0_r71_c33;
    wire stage0_r65_c40;
    wire stage0_r66_c39;
    wire stage0_r67_c38;
    wire stage0_r68_c37;
    wire stage0_r69_c36;
    wire stage0_r70_c35;
    wire stage0_r71_c34;
    wire stage0_r66_c40;
    wire stage0_r67_c39;
    wire stage0_r68_c38;
    wire stage0_r69_c37;
    wire stage0_r70_c36;
    wire stage0_r71_c35;
    wire stage0_r67_c40;
    wire stage0_r68_c39;
    wire stage0_r69_c38;
    wire stage0_r70_c37;
    wire stage0_r71_c36;
    wire stage0_r68_c40;
    wire stage0_r69_c39;
    wire stage0_r70_c38;
    wire stage0_r71_c37;
    wire stage0_r69_c40;
    wire stage0_r70_c39;
    wire stage0_r71_c38;
    wire stage0_r70_c40;
    wire stage0_r71_c39;
    wire stage0_r71_c40;
    wire stage1_c1_s_ha0;
    wire stage1_c1_c_ha0;
    wire stage1_c2_s_fa0;
    wire stage1_c2_c_fa0;
    wire stage1_c3_s_fa0;
    wire stage1_c3_c_fa0;
    wire stage1_c4_s_fa0;
    wire stage1_c4_c_fa0;
    wire stage1_c4_s_ha0;
    wire stage1_c4_c_ha0;
    wire stage1_c5_s_fa0;
    wire stage1_c5_c_fa0;
    wire stage1_c5_s_fa1;
    wire stage1_c5_c_fa1;
    wire stage1_c6_s_fa0;
    wire stage1_c6_c_fa0;
    wire stage1_c6_s_fa1;
    wire stage1_c6_c_fa1;
    wire stage1_c7_s_fa0;
    wire stage1_c7_c_fa0;
    wire stage1_c7_s_fa1;
    wire stage1_c7_c_fa1;
    wire stage1_c7_s_ha0;
    wire stage1_c7_c_ha0;
    wire stage1_c8_s_fa0;
    wire stage1_c8_c_fa0;
    wire stage1_c8_s_fa1;
    wire stage1_c8_c_fa1;
    wire stage1_c8_s_fa2;
    wire stage1_c8_c_fa2;
    wire stage1_c9_s_fa0;
    wire stage1_c9_c_fa0;
    wire stage1_c9_s_fa1;
    wire stage1_c9_c_fa1;
    wire stage1_c9_s_fa2;
    wire stage1_c9_c_fa2;
    wire stage1_c10_s_fa0;
    wire stage1_c10_c_fa0;
    wire stage1_c10_s_fa1;
    wire stage1_c10_c_fa1;
    wire stage1_c10_s_fa2;
    wire stage1_c10_c_fa2;
    wire stage1_c10_s_ha0;
    wire stage1_c10_c_ha0;
    wire stage1_c11_s_fa0;
    wire stage1_c11_c_fa0;
    wire stage1_c11_s_fa1;
    wire stage1_c11_c_fa1;
    wire stage1_c11_s_fa2;
    wire stage1_c11_c_fa2;
    wire stage1_c11_s_fa3;
    wire stage1_c11_c_fa3;
    wire stage1_c12_s_fa0;
    wire stage1_c12_c_fa0;
    wire stage1_c12_s_fa1;
    wire stage1_c12_c_fa1;
    wire stage1_c12_s_fa2;
    wire stage1_c12_c_fa2;
    wire stage1_c12_s_fa3;
    wire stage1_c12_c_fa3;
    wire stage1_c13_s_fa0;
    wire stage1_c13_c_fa0;
    wire stage1_c13_s_fa1;
    wire stage1_c13_c_fa1;
    wire stage1_c13_s_fa2;
    wire stage1_c13_c_fa2;
    wire stage1_c13_s_fa3;
    wire stage1_c13_c_fa3;
    wire stage1_c13_s_ha0;
    wire stage1_c13_c_ha0;
    wire stage1_c14_s_fa0;
    wire stage1_c14_c_fa0;
    wire stage1_c14_s_fa1;
    wire stage1_c14_c_fa1;
    wire stage1_c14_s_fa2;
    wire stage1_c14_c_fa2;
    wire stage1_c14_s_fa3;
    wire stage1_c14_c_fa3;
    wire stage1_c14_s_fa4;
    wire stage1_c14_c_fa4;
    wire stage1_c15_s_fa0;
    wire stage1_c15_c_fa0;
    wire stage1_c15_s_fa1;
    wire stage1_c15_c_fa1;
    wire stage1_c15_s_fa2;
    wire stage1_c15_c_fa2;
    wire stage1_c15_s_fa3;
    wire stage1_c15_c_fa3;
    wire stage1_c15_s_fa4;
    wire stage1_c15_c_fa4;
    wire stage1_c16_s_fa0;
    wire stage1_c16_c_fa0;
    wire stage1_c16_s_fa1;
    wire stage1_c16_c_fa1;
    wire stage1_c16_s_fa2;
    wire stage1_c16_c_fa2;
    wire stage1_c16_s_fa3;
    wire stage1_c16_c_fa3;
    wire stage1_c16_s_fa4;
    wire stage1_c16_c_fa4;
    wire stage1_c16_s_ha0;
    wire stage1_c16_c_ha0;
    wire stage1_c17_s_fa0;
    wire stage1_c17_c_fa0;
    wire stage1_c17_s_fa1;
    wire stage1_c17_c_fa1;
    wire stage1_c17_s_fa2;
    wire stage1_c17_c_fa2;
    wire stage1_c17_s_fa3;
    wire stage1_c17_c_fa3;
    wire stage1_c17_s_fa4;
    wire stage1_c17_c_fa4;
    wire stage1_c17_s_fa5;
    wire stage1_c17_c_fa5;
    wire stage1_c18_s_fa0;
    wire stage1_c18_c_fa0;
    wire stage1_c18_s_fa1;
    wire stage1_c18_c_fa1;
    wire stage1_c18_s_fa2;
    wire stage1_c18_c_fa2;
    wire stage1_c18_s_fa3;
    wire stage1_c18_c_fa3;
    wire stage1_c18_s_fa4;
    wire stage1_c18_c_fa4;
    wire stage1_c18_s_fa5;
    wire stage1_c18_c_fa5;
    wire stage1_c19_s_fa0;
    wire stage1_c19_c_fa0;
    wire stage1_c19_s_fa1;
    wire stage1_c19_c_fa1;
    wire stage1_c19_s_fa2;
    wire stage1_c19_c_fa2;
    wire stage1_c19_s_fa3;
    wire stage1_c19_c_fa3;
    wire stage1_c19_s_fa4;
    wire stage1_c19_c_fa4;
    wire stage1_c19_s_fa5;
    wire stage1_c19_c_fa5;
    wire stage1_c19_s_ha0;
    wire stage1_c19_c_ha0;
    wire stage1_c20_s_fa0;
    wire stage1_c20_c_fa0;
    wire stage1_c20_s_fa1;
    wire stage1_c20_c_fa1;
    wire stage1_c20_s_fa2;
    wire stage1_c20_c_fa2;
    wire stage1_c20_s_fa3;
    wire stage1_c20_c_fa3;
    wire stage1_c20_s_fa4;
    wire stage1_c20_c_fa4;
    wire stage1_c20_s_fa5;
    wire stage1_c20_c_fa5;
    wire stage1_c20_s_fa6;
    wire stage1_c20_c_fa6;
    wire stage1_c21_s_fa0;
    wire stage1_c21_c_fa0;
    wire stage1_c21_s_fa1;
    wire stage1_c21_c_fa1;
    wire stage1_c21_s_fa2;
    wire stage1_c21_c_fa2;
    wire stage1_c21_s_fa3;
    wire stage1_c21_c_fa3;
    wire stage1_c21_s_fa4;
    wire stage1_c21_c_fa4;
    wire stage1_c21_s_fa5;
    wire stage1_c21_c_fa5;
    wire stage1_c21_s_fa6;
    wire stage1_c21_c_fa6;
    wire stage1_c22_s_fa0;
    wire stage1_c22_c_fa0;
    wire stage1_c22_s_fa1;
    wire stage1_c22_c_fa1;
    wire stage1_c22_s_fa2;
    wire stage1_c22_c_fa2;
    wire stage1_c22_s_fa3;
    wire stage1_c22_c_fa3;
    wire stage1_c22_s_fa4;
    wire stage1_c22_c_fa4;
    wire stage1_c22_s_fa5;
    wire stage1_c22_c_fa5;
    wire stage1_c22_s_fa6;
    wire stage1_c22_c_fa6;
    wire stage1_c22_s_ha0;
    wire stage1_c22_c_ha0;
    wire stage1_c23_s_fa0;
    wire stage1_c23_c_fa0;
    wire stage1_c23_s_fa1;
    wire stage1_c23_c_fa1;
    wire stage1_c23_s_fa2;
    wire stage1_c23_c_fa2;
    wire stage1_c23_s_fa3;
    wire stage1_c23_c_fa3;
    wire stage1_c23_s_fa4;
    wire stage1_c23_c_fa4;
    wire stage1_c23_s_fa5;
    wire stage1_c23_c_fa5;
    wire stage1_c23_s_fa6;
    wire stage1_c23_c_fa6;
    wire stage1_c23_s_fa7;
    wire stage1_c23_c_fa7;
    wire stage1_c24_s_fa0;
    wire stage1_c24_c_fa0;
    wire stage1_c24_s_fa1;
    wire stage1_c24_c_fa1;
    wire stage1_c24_s_fa2;
    wire stage1_c24_c_fa2;
    wire stage1_c24_s_fa3;
    wire stage1_c24_c_fa3;
    wire stage1_c24_s_fa4;
    wire stage1_c24_c_fa4;
    wire stage1_c24_s_fa5;
    wire stage1_c24_c_fa5;
    wire stage1_c24_s_fa6;
    wire stage1_c24_c_fa6;
    wire stage1_c24_s_fa7;
    wire stage1_c24_c_fa7;
    wire stage1_c25_s_fa0;
    wire stage1_c25_c_fa0;
    wire stage1_c25_s_fa1;
    wire stage1_c25_c_fa1;
    wire stage1_c25_s_fa2;
    wire stage1_c25_c_fa2;
    wire stage1_c25_s_fa3;
    wire stage1_c25_c_fa3;
    wire stage1_c25_s_fa4;
    wire stage1_c25_c_fa4;
    wire stage1_c25_s_fa5;
    wire stage1_c25_c_fa5;
    wire stage1_c25_s_fa6;
    wire stage1_c25_c_fa6;
    wire stage1_c25_s_fa7;
    wire stage1_c25_c_fa7;
    wire stage1_c25_s_ha0;
    wire stage1_c25_c_ha0;
    wire stage1_c26_s_fa0;
    wire stage1_c26_c_fa0;
    wire stage1_c26_s_fa1;
    wire stage1_c26_c_fa1;
    wire stage1_c26_s_fa2;
    wire stage1_c26_c_fa2;
    wire stage1_c26_s_fa3;
    wire stage1_c26_c_fa3;
    wire stage1_c26_s_fa4;
    wire stage1_c26_c_fa4;
    wire stage1_c26_s_fa5;
    wire stage1_c26_c_fa5;
    wire stage1_c26_s_fa6;
    wire stage1_c26_c_fa6;
    wire stage1_c26_s_fa7;
    wire stage1_c26_c_fa7;
    wire stage1_c26_s_fa8;
    wire stage1_c26_c_fa8;
    wire stage1_c27_s_fa0;
    wire stage1_c27_c_fa0;
    wire stage1_c27_s_fa1;
    wire stage1_c27_c_fa1;
    wire stage1_c27_s_fa2;
    wire stage1_c27_c_fa2;
    wire stage1_c27_s_fa3;
    wire stage1_c27_c_fa3;
    wire stage1_c27_s_fa4;
    wire stage1_c27_c_fa4;
    wire stage1_c27_s_fa5;
    wire stage1_c27_c_fa5;
    wire stage1_c27_s_fa6;
    wire stage1_c27_c_fa6;
    wire stage1_c27_s_fa7;
    wire stage1_c27_c_fa7;
    wire stage1_c27_s_fa8;
    wire stage1_c27_c_fa8;
    wire stage1_c28_s_fa0;
    wire stage1_c28_c_fa0;
    wire stage1_c28_s_fa1;
    wire stage1_c28_c_fa1;
    wire stage1_c28_s_fa2;
    wire stage1_c28_c_fa2;
    wire stage1_c28_s_fa3;
    wire stage1_c28_c_fa3;
    wire stage1_c28_s_fa4;
    wire stage1_c28_c_fa4;
    wire stage1_c28_s_fa5;
    wire stage1_c28_c_fa5;
    wire stage1_c28_s_fa6;
    wire stage1_c28_c_fa6;
    wire stage1_c28_s_fa7;
    wire stage1_c28_c_fa7;
    wire stage1_c28_s_fa8;
    wire stage1_c28_c_fa8;
    wire stage1_c28_s_ha0;
    wire stage1_c28_c_ha0;
    wire stage1_c29_s_fa0;
    wire stage1_c29_c_fa0;
    wire stage1_c29_s_fa1;
    wire stage1_c29_c_fa1;
    wire stage1_c29_s_fa2;
    wire stage1_c29_c_fa2;
    wire stage1_c29_s_fa3;
    wire stage1_c29_c_fa3;
    wire stage1_c29_s_fa4;
    wire stage1_c29_c_fa4;
    wire stage1_c29_s_fa5;
    wire stage1_c29_c_fa5;
    wire stage1_c29_s_fa6;
    wire stage1_c29_c_fa6;
    wire stage1_c29_s_fa7;
    wire stage1_c29_c_fa7;
    wire stage1_c29_s_fa8;
    wire stage1_c29_c_fa8;
    wire stage1_c29_s_fa9;
    wire stage1_c29_c_fa9;
    wire stage1_c30_s_fa0;
    wire stage1_c30_c_fa0;
    wire stage1_c30_s_fa1;
    wire stage1_c30_c_fa1;
    wire stage1_c30_s_fa2;
    wire stage1_c30_c_fa2;
    wire stage1_c30_s_fa3;
    wire stage1_c30_c_fa3;
    wire stage1_c30_s_fa4;
    wire stage1_c30_c_fa4;
    wire stage1_c30_s_fa5;
    wire stage1_c30_c_fa5;
    wire stage1_c30_s_fa6;
    wire stage1_c30_c_fa6;
    wire stage1_c30_s_fa7;
    wire stage1_c30_c_fa7;
    wire stage1_c30_s_fa8;
    wire stage1_c30_c_fa8;
    wire stage1_c30_s_fa9;
    wire stage1_c30_c_fa9;
    wire stage1_c31_s_fa0;
    wire stage1_c31_c_fa0;
    wire stage1_c31_s_fa1;
    wire stage1_c31_c_fa1;
    wire stage1_c31_s_fa2;
    wire stage1_c31_c_fa2;
    wire stage1_c31_s_fa3;
    wire stage1_c31_c_fa3;
    wire stage1_c31_s_fa4;
    wire stage1_c31_c_fa4;
    wire stage1_c31_s_fa5;
    wire stage1_c31_c_fa5;
    wire stage1_c31_s_fa6;
    wire stage1_c31_c_fa6;
    wire stage1_c31_s_fa7;
    wire stage1_c31_c_fa7;
    wire stage1_c31_s_fa8;
    wire stage1_c31_c_fa8;
    wire stage1_c31_s_fa9;
    wire stage1_c31_c_fa9;
    wire stage1_c31_s_ha0;
    wire stage1_c31_c_ha0;
    wire stage1_c32_s_fa0;
    wire stage1_c32_c_fa0;
    wire stage1_c32_s_fa1;
    wire stage1_c32_c_fa1;
    wire stage1_c32_s_fa2;
    wire stage1_c32_c_fa2;
    wire stage1_c32_s_fa3;
    wire stage1_c32_c_fa3;
    wire stage1_c32_s_fa4;
    wire stage1_c32_c_fa4;
    wire stage1_c32_s_fa5;
    wire stage1_c32_c_fa5;
    wire stage1_c32_s_fa6;
    wire stage1_c32_c_fa6;
    wire stage1_c32_s_fa7;
    wire stage1_c32_c_fa7;
    wire stage1_c32_s_fa8;
    wire stage1_c32_c_fa8;
    wire stage1_c32_s_fa9;
    wire stage1_c32_c_fa9;
    wire stage1_c32_s_fa10;
    wire stage1_c32_c_fa10;
    wire stage1_c33_s_fa0;
    wire stage1_c33_c_fa0;
    wire stage1_c33_s_fa1;
    wire stage1_c33_c_fa1;
    wire stage1_c33_s_fa2;
    wire stage1_c33_c_fa2;
    wire stage1_c33_s_fa3;
    wire stage1_c33_c_fa3;
    wire stage1_c33_s_fa4;
    wire stage1_c33_c_fa4;
    wire stage1_c33_s_fa5;
    wire stage1_c33_c_fa5;
    wire stage1_c33_s_fa6;
    wire stage1_c33_c_fa6;
    wire stage1_c33_s_fa7;
    wire stage1_c33_c_fa7;
    wire stage1_c33_s_fa8;
    wire stage1_c33_c_fa8;
    wire stage1_c33_s_fa9;
    wire stage1_c33_c_fa9;
    wire stage1_c33_s_fa10;
    wire stage1_c33_c_fa10;
    wire stage1_c34_s_fa0;
    wire stage1_c34_c_fa0;
    wire stage1_c34_s_fa1;
    wire stage1_c34_c_fa1;
    wire stage1_c34_s_fa2;
    wire stage1_c34_c_fa2;
    wire stage1_c34_s_fa3;
    wire stage1_c34_c_fa3;
    wire stage1_c34_s_fa4;
    wire stage1_c34_c_fa4;
    wire stage1_c34_s_fa5;
    wire stage1_c34_c_fa5;
    wire stage1_c34_s_fa6;
    wire stage1_c34_c_fa6;
    wire stage1_c34_s_fa7;
    wire stage1_c34_c_fa7;
    wire stage1_c34_s_fa8;
    wire stage1_c34_c_fa8;
    wire stage1_c34_s_fa9;
    wire stage1_c34_c_fa9;
    wire stage1_c34_s_fa10;
    wire stage1_c34_c_fa10;
    wire stage1_c34_s_ha0;
    wire stage1_c34_c_ha0;
    wire stage1_c35_s_fa0;
    wire stage1_c35_c_fa0;
    wire stage1_c35_s_fa1;
    wire stage1_c35_c_fa1;
    wire stage1_c35_s_fa2;
    wire stage1_c35_c_fa2;
    wire stage1_c35_s_fa3;
    wire stage1_c35_c_fa3;
    wire stage1_c35_s_fa4;
    wire stage1_c35_c_fa4;
    wire stage1_c35_s_fa5;
    wire stage1_c35_c_fa5;
    wire stage1_c35_s_fa6;
    wire stage1_c35_c_fa6;
    wire stage1_c35_s_fa7;
    wire stage1_c35_c_fa7;
    wire stage1_c35_s_fa8;
    wire stage1_c35_c_fa8;
    wire stage1_c35_s_fa9;
    wire stage1_c35_c_fa9;
    wire stage1_c35_s_fa10;
    wire stage1_c35_c_fa10;
    wire stage1_c35_s_fa11;
    wire stage1_c35_c_fa11;
    wire stage1_c36_s_fa0;
    wire stage1_c36_c_fa0;
    wire stage1_c36_s_fa1;
    wire stage1_c36_c_fa1;
    wire stage1_c36_s_fa2;
    wire stage1_c36_c_fa2;
    wire stage1_c36_s_fa3;
    wire stage1_c36_c_fa3;
    wire stage1_c36_s_fa4;
    wire stage1_c36_c_fa4;
    wire stage1_c36_s_fa5;
    wire stage1_c36_c_fa5;
    wire stage1_c36_s_fa6;
    wire stage1_c36_c_fa6;
    wire stage1_c36_s_fa7;
    wire stage1_c36_c_fa7;
    wire stage1_c36_s_fa8;
    wire stage1_c36_c_fa8;
    wire stage1_c36_s_fa9;
    wire stage1_c36_c_fa9;
    wire stage1_c36_s_fa10;
    wire stage1_c36_c_fa10;
    wire stage1_c36_s_fa11;
    wire stage1_c36_c_fa11;
    wire stage1_c37_s_fa0;
    wire stage1_c37_c_fa0;
    wire stage1_c37_s_fa1;
    wire stage1_c37_c_fa1;
    wire stage1_c37_s_fa2;
    wire stage1_c37_c_fa2;
    wire stage1_c37_s_fa3;
    wire stage1_c37_c_fa3;
    wire stage1_c37_s_fa4;
    wire stage1_c37_c_fa4;
    wire stage1_c37_s_fa5;
    wire stage1_c37_c_fa5;
    wire stage1_c37_s_fa6;
    wire stage1_c37_c_fa6;
    wire stage1_c37_s_fa7;
    wire stage1_c37_c_fa7;
    wire stage1_c37_s_fa8;
    wire stage1_c37_c_fa8;
    wire stage1_c37_s_fa9;
    wire stage1_c37_c_fa9;
    wire stage1_c37_s_fa10;
    wire stage1_c37_c_fa10;
    wire stage1_c37_s_fa11;
    wire stage1_c37_c_fa11;
    wire stage1_c37_s_ha0;
    wire stage1_c37_c_ha0;
    wire stage1_c38_s_fa0;
    wire stage1_c38_c_fa0;
    wire stage1_c38_s_fa1;
    wire stage1_c38_c_fa1;
    wire stage1_c38_s_fa2;
    wire stage1_c38_c_fa2;
    wire stage1_c38_s_fa3;
    wire stage1_c38_c_fa3;
    wire stage1_c38_s_fa4;
    wire stage1_c38_c_fa4;
    wire stage1_c38_s_fa5;
    wire stage1_c38_c_fa5;
    wire stage1_c38_s_fa6;
    wire stage1_c38_c_fa6;
    wire stage1_c38_s_fa7;
    wire stage1_c38_c_fa7;
    wire stage1_c38_s_fa8;
    wire stage1_c38_c_fa8;
    wire stage1_c38_s_fa9;
    wire stage1_c38_c_fa9;
    wire stage1_c38_s_fa10;
    wire stage1_c38_c_fa10;
    wire stage1_c38_s_fa11;
    wire stage1_c38_c_fa11;
    wire stage1_c38_s_fa12;
    wire stage1_c38_c_fa12;
    wire stage1_c39_s_fa0;
    wire stage1_c39_c_fa0;
    wire stage1_c39_s_fa1;
    wire stage1_c39_c_fa1;
    wire stage1_c39_s_fa2;
    wire stage1_c39_c_fa2;
    wire stage1_c39_s_fa3;
    wire stage1_c39_c_fa3;
    wire stage1_c39_s_fa4;
    wire stage1_c39_c_fa4;
    wire stage1_c39_s_fa5;
    wire stage1_c39_c_fa5;
    wire stage1_c39_s_fa6;
    wire stage1_c39_c_fa6;
    wire stage1_c39_s_fa7;
    wire stage1_c39_c_fa7;
    wire stage1_c39_s_fa8;
    wire stage1_c39_c_fa8;
    wire stage1_c39_s_fa9;
    wire stage1_c39_c_fa9;
    wire stage1_c39_s_fa10;
    wire stage1_c39_c_fa10;
    wire stage1_c39_s_fa11;
    wire stage1_c39_c_fa11;
    wire stage1_c39_s_fa12;
    wire stage1_c39_c_fa12;
    wire stage1_c40_s_fa0;
    wire stage1_c40_c_fa0;
    wire stage1_c40_s_fa1;
    wire stage1_c40_c_fa1;
    wire stage1_c40_s_fa2;
    wire stage1_c40_c_fa2;
    wire stage1_c40_s_fa3;
    wire stage1_c40_c_fa3;
    wire stage1_c40_s_fa4;
    wire stage1_c40_c_fa4;
    wire stage1_c40_s_fa5;
    wire stage1_c40_c_fa5;
    wire stage1_c40_s_fa6;
    wire stage1_c40_c_fa6;
    wire stage1_c40_s_fa7;
    wire stage1_c40_c_fa7;
    wire stage1_c40_s_fa8;
    wire stage1_c40_c_fa8;
    wire stage1_c40_s_fa9;
    wire stage1_c40_c_fa9;
    wire stage1_c40_s_fa10;
    wire stage1_c40_c_fa10;
    wire stage1_c40_s_fa11;
    wire stage1_c40_c_fa11;
    wire stage1_c40_s_fa12;
    wire stage1_c40_c_fa12;
    wire stage1_c40_s_ha0;
    wire stage1_c40_c_ha0;
    wire stage1_c41_s_fa0;
    wire stage1_c41_c_fa0;
    wire stage1_c41_s_fa1;
    wire stage1_c41_c_fa1;
    wire stage1_c41_s_fa2;
    wire stage1_c41_c_fa2;
    wire stage1_c41_s_fa3;
    wire stage1_c41_c_fa3;
    wire stage1_c41_s_fa4;
    wire stage1_c41_c_fa4;
    wire stage1_c41_s_fa5;
    wire stage1_c41_c_fa5;
    wire stage1_c41_s_fa6;
    wire stage1_c41_c_fa6;
    wire stage1_c41_s_fa7;
    wire stage1_c41_c_fa7;
    wire stage1_c41_s_fa8;
    wire stage1_c41_c_fa8;
    wire stage1_c41_s_fa9;
    wire stage1_c41_c_fa9;
    wire stage1_c41_s_fa10;
    wire stage1_c41_c_fa10;
    wire stage1_c41_s_fa11;
    wire stage1_c41_c_fa11;
    wire stage1_c41_s_fa12;
    wire stage1_c41_c_fa12;
    wire stage1_c41_s_ha0;
    wire stage1_c41_c_ha0;
    wire stage1_c42_s_fa0;
    wire stage1_c42_c_fa0;
    wire stage1_c42_s_fa1;
    wire stage1_c42_c_fa1;
    wire stage1_c42_s_fa2;
    wire stage1_c42_c_fa2;
    wire stage1_c42_s_fa3;
    wire stage1_c42_c_fa3;
    wire stage1_c42_s_fa4;
    wire stage1_c42_c_fa4;
    wire stage1_c42_s_fa5;
    wire stage1_c42_c_fa5;
    wire stage1_c42_s_fa6;
    wire stage1_c42_c_fa6;
    wire stage1_c42_s_fa7;
    wire stage1_c42_c_fa7;
    wire stage1_c42_s_fa8;
    wire stage1_c42_c_fa8;
    wire stage1_c42_s_fa9;
    wire stage1_c42_c_fa9;
    wire stage1_c42_s_fa10;
    wire stage1_c42_c_fa10;
    wire stage1_c42_s_fa11;
    wire stage1_c42_c_fa11;
    wire stage1_c42_s_fa12;
    wire stage1_c42_c_fa12;
    wire stage1_c42_s_ha0;
    wire stage1_c42_c_ha0;
    wire stage1_c43_s_fa0;
    wire stage1_c43_c_fa0;
    wire stage1_c43_s_fa1;
    wire stage1_c43_c_fa1;
    wire stage1_c43_s_fa2;
    wire stage1_c43_c_fa2;
    wire stage1_c43_s_fa3;
    wire stage1_c43_c_fa3;
    wire stage1_c43_s_fa4;
    wire stage1_c43_c_fa4;
    wire stage1_c43_s_fa5;
    wire stage1_c43_c_fa5;
    wire stage1_c43_s_fa6;
    wire stage1_c43_c_fa6;
    wire stage1_c43_s_fa7;
    wire stage1_c43_c_fa7;
    wire stage1_c43_s_fa8;
    wire stage1_c43_c_fa8;
    wire stage1_c43_s_fa9;
    wire stage1_c43_c_fa9;
    wire stage1_c43_s_fa10;
    wire stage1_c43_c_fa10;
    wire stage1_c43_s_fa11;
    wire stage1_c43_c_fa11;
    wire stage1_c43_s_fa12;
    wire stage1_c43_c_fa12;
    wire stage1_c43_s_ha0;
    wire stage1_c43_c_ha0;
    wire stage1_c44_s_fa0;
    wire stage1_c44_c_fa0;
    wire stage1_c44_s_fa1;
    wire stage1_c44_c_fa1;
    wire stage1_c44_s_fa2;
    wire stage1_c44_c_fa2;
    wire stage1_c44_s_fa3;
    wire stage1_c44_c_fa3;
    wire stage1_c44_s_fa4;
    wire stage1_c44_c_fa4;
    wire stage1_c44_s_fa5;
    wire stage1_c44_c_fa5;
    wire stage1_c44_s_fa6;
    wire stage1_c44_c_fa6;
    wire stage1_c44_s_fa7;
    wire stage1_c44_c_fa7;
    wire stage1_c44_s_fa8;
    wire stage1_c44_c_fa8;
    wire stage1_c44_s_fa9;
    wire stage1_c44_c_fa9;
    wire stage1_c44_s_fa10;
    wire stage1_c44_c_fa10;
    wire stage1_c44_s_fa11;
    wire stage1_c44_c_fa11;
    wire stage1_c44_s_fa12;
    wire stage1_c44_c_fa12;
    wire stage1_c44_s_ha0;
    wire stage1_c44_c_ha0;
    wire stage1_c45_s_fa0;
    wire stage1_c45_c_fa0;
    wire stage1_c45_s_fa1;
    wire stage1_c45_c_fa1;
    wire stage1_c45_s_fa2;
    wire stage1_c45_c_fa2;
    wire stage1_c45_s_fa3;
    wire stage1_c45_c_fa3;
    wire stage1_c45_s_fa4;
    wire stage1_c45_c_fa4;
    wire stage1_c45_s_fa5;
    wire stage1_c45_c_fa5;
    wire stage1_c45_s_fa6;
    wire stage1_c45_c_fa6;
    wire stage1_c45_s_fa7;
    wire stage1_c45_c_fa7;
    wire stage1_c45_s_fa8;
    wire stage1_c45_c_fa8;
    wire stage1_c45_s_fa9;
    wire stage1_c45_c_fa9;
    wire stage1_c45_s_fa10;
    wire stage1_c45_c_fa10;
    wire stage1_c45_s_fa11;
    wire stage1_c45_c_fa11;
    wire stage1_c45_s_fa12;
    wire stage1_c45_c_fa12;
    wire stage1_c45_s_ha0;
    wire stage1_c45_c_ha0;
    wire stage1_c46_s_fa0;
    wire stage1_c46_c_fa0;
    wire stage1_c46_s_fa1;
    wire stage1_c46_c_fa1;
    wire stage1_c46_s_fa2;
    wire stage1_c46_c_fa2;
    wire stage1_c46_s_fa3;
    wire stage1_c46_c_fa3;
    wire stage1_c46_s_fa4;
    wire stage1_c46_c_fa4;
    wire stage1_c46_s_fa5;
    wire stage1_c46_c_fa5;
    wire stage1_c46_s_fa6;
    wire stage1_c46_c_fa6;
    wire stage1_c46_s_fa7;
    wire stage1_c46_c_fa7;
    wire stage1_c46_s_fa8;
    wire stage1_c46_c_fa8;
    wire stage1_c46_s_fa9;
    wire stage1_c46_c_fa9;
    wire stage1_c46_s_fa10;
    wire stage1_c46_c_fa10;
    wire stage1_c46_s_fa11;
    wire stage1_c46_c_fa11;
    wire stage1_c46_s_fa12;
    wire stage1_c46_c_fa12;
    wire stage1_c46_s_ha0;
    wire stage1_c46_c_ha0;
    wire stage1_c47_s_fa0;
    wire stage1_c47_c_fa0;
    wire stage1_c47_s_fa1;
    wire stage1_c47_c_fa1;
    wire stage1_c47_s_fa2;
    wire stage1_c47_c_fa2;
    wire stage1_c47_s_fa3;
    wire stage1_c47_c_fa3;
    wire stage1_c47_s_fa4;
    wire stage1_c47_c_fa4;
    wire stage1_c47_s_fa5;
    wire stage1_c47_c_fa5;
    wire stage1_c47_s_fa6;
    wire stage1_c47_c_fa6;
    wire stage1_c47_s_fa7;
    wire stage1_c47_c_fa7;
    wire stage1_c47_s_fa8;
    wire stage1_c47_c_fa8;
    wire stage1_c47_s_fa9;
    wire stage1_c47_c_fa9;
    wire stage1_c47_s_fa10;
    wire stage1_c47_c_fa10;
    wire stage1_c47_s_fa11;
    wire stage1_c47_c_fa11;
    wire stage1_c47_s_fa12;
    wire stage1_c47_c_fa12;
    wire stage1_c47_s_ha0;
    wire stage1_c47_c_ha0;
    wire stage1_c48_s_fa0;
    wire stage1_c48_c_fa0;
    wire stage1_c48_s_fa1;
    wire stage1_c48_c_fa1;
    wire stage1_c48_s_fa2;
    wire stage1_c48_c_fa2;
    wire stage1_c48_s_fa3;
    wire stage1_c48_c_fa3;
    wire stage1_c48_s_fa4;
    wire stage1_c48_c_fa4;
    wire stage1_c48_s_fa5;
    wire stage1_c48_c_fa5;
    wire stage1_c48_s_fa6;
    wire stage1_c48_c_fa6;
    wire stage1_c48_s_fa7;
    wire stage1_c48_c_fa7;
    wire stage1_c48_s_fa8;
    wire stage1_c48_c_fa8;
    wire stage1_c48_s_fa9;
    wire stage1_c48_c_fa9;
    wire stage1_c48_s_fa10;
    wire stage1_c48_c_fa10;
    wire stage1_c48_s_fa11;
    wire stage1_c48_c_fa11;
    wire stage1_c48_s_fa12;
    wire stage1_c48_c_fa12;
    wire stage1_c48_s_ha0;
    wire stage1_c48_c_ha0;
    wire stage1_c49_s_fa0;
    wire stage1_c49_c_fa0;
    wire stage1_c49_s_fa1;
    wire stage1_c49_c_fa1;
    wire stage1_c49_s_fa2;
    wire stage1_c49_c_fa2;
    wire stage1_c49_s_fa3;
    wire stage1_c49_c_fa3;
    wire stage1_c49_s_fa4;
    wire stage1_c49_c_fa4;
    wire stage1_c49_s_fa5;
    wire stage1_c49_c_fa5;
    wire stage1_c49_s_fa6;
    wire stage1_c49_c_fa6;
    wire stage1_c49_s_fa7;
    wire stage1_c49_c_fa7;
    wire stage1_c49_s_fa8;
    wire stage1_c49_c_fa8;
    wire stage1_c49_s_fa9;
    wire stage1_c49_c_fa9;
    wire stage1_c49_s_fa10;
    wire stage1_c49_c_fa10;
    wire stage1_c49_s_fa11;
    wire stage1_c49_c_fa11;
    wire stage1_c49_s_fa12;
    wire stage1_c49_c_fa12;
    wire stage1_c49_s_ha0;
    wire stage1_c49_c_ha0;
    wire stage1_c50_s_fa0;
    wire stage1_c50_c_fa0;
    wire stage1_c50_s_fa1;
    wire stage1_c50_c_fa1;
    wire stage1_c50_s_fa2;
    wire stage1_c50_c_fa2;
    wire stage1_c50_s_fa3;
    wire stage1_c50_c_fa3;
    wire stage1_c50_s_fa4;
    wire stage1_c50_c_fa4;
    wire stage1_c50_s_fa5;
    wire stage1_c50_c_fa5;
    wire stage1_c50_s_fa6;
    wire stage1_c50_c_fa6;
    wire stage1_c50_s_fa7;
    wire stage1_c50_c_fa7;
    wire stage1_c50_s_fa8;
    wire stage1_c50_c_fa8;
    wire stage1_c50_s_fa9;
    wire stage1_c50_c_fa9;
    wire stage1_c50_s_fa10;
    wire stage1_c50_c_fa10;
    wire stage1_c50_s_fa11;
    wire stage1_c50_c_fa11;
    wire stage1_c50_s_fa12;
    wire stage1_c50_c_fa12;
    wire stage1_c50_s_ha0;
    wire stage1_c50_c_ha0;
    wire stage1_c51_s_fa0;
    wire stage1_c51_c_fa0;
    wire stage1_c51_s_fa1;
    wire stage1_c51_c_fa1;
    wire stage1_c51_s_fa2;
    wire stage1_c51_c_fa2;
    wire stage1_c51_s_fa3;
    wire stage1_c51_c_fa3;
    wire stage1_c51_s_fa4;
    wire stage1_c51_c_fa4;
    wire stage1_c51_s_fa5;
    wire stage1_c51_c_fa5;
    wire stage1_c51_s_fa6;
    wire stage1_c51_c_fa6;
    wire stage1_c51_s_fa7;
    wire stage1_c51_c_fa7;
    wire stage1_c51_s_fa8;
    wire stage1_c51_c_fa8;
    wire stage1_c51_s_fa9;
    wire stage1_c51_c_fa9;
    wire stage1_c51_s_fa10;
    wire stage1_c51_c_fa10;
    wire stage1_c51_s_fa11;
    wire stage1_c51_c_fa11;
    wire stage1_c51_s_fa12;
    wire stage1_c51_c_fa12;
    wire stage1_c51_s_ha0;
    wire stage1_c51_c_ha0;
    wire stage1_c52_s_fa0;
    wire stage1_c52_c_fa0;
    wire stage1_c52_s_fa1;
    wire stage1_c52_c_fa1;
    wire stage1_c52_s_fa2;
    wire stage1_c52_c_fa2;
    wire stage1_c52_s_fa3;
    wire stage1_c52_c_fa3;
    wire stage1_c52_s_fa4;
    wire stage1_c52_c_fa4;
    wire stage1_c52_s_fa5;
    wire stage1_c52_c_fa5;
    wire stage1_c52_s_fa6;
    wire stage1_c52_c_fa6;
    wire stage1_c52_s_fa7;
    wire stage1_c52_c_fa7;
    wire stage1_c52_s_fa8;
    wire stage1_c52_c_fa8;
    wire stage1_c52_s_fa9;
    wire stage1_c52_c_fa9;
    wire stage1_c52_s_fa10;
    wire stage1_c52_c_fa10;
    wire stage1_c52_s_fa11;
    wire stage1_c52_c_fa11;
    wire stage1_c52_s_fa12;
    wire stage1_c52_c_fa12;
    wire stage1_c52_s_ha0;
    wire stage1_c52_c_ha0;
    wire stage1_c53_s_fa0;
    wire stage1_c53_c_fa0;
    wire stage1_c53_s_fa1;
    wire stage1_c53_c_fa1;
    wire stage1_c53_s_fa2;
    wire stage1_c53_c_fa2;
    wire stage1_c53_s_fa3;
    wire stage1_c53_c_fa3;
    wire stage1_c53_s_fa4;
    wire stage1_c53_c_fa4;
    wire stage1_c53_s_fa5;
    wire stage1_c53_c_fa5;
    wire stage1_c53_s_fa6;
    wire stage1_c53_c_fa6;
    wire stage1_c53_s_fa7;
    wire stage1_c53_c_fa7;
    wire stage1_c53_s_fa8;
    wire stage1_c53_c_fa8;
    wire stage1_c53_s_fa9;
    wire stage1_c53_c_fa9;
    wire stage1_c53_s_fa10;
    wire stage1_c53_c_fa10;
    wire stage1_c53_s_fa11;
    wire stage1_c53_c_fa11;
    wire stage1_c53_s_fa12;
    wire stage1_c53_c_fa12;
    wire stage1_c53_s_ha0;
    wire stage1_c53_c_ha0;
    wire stage1_c54_s_fa0;
    wire stage1_c54_c_fa0;
    wire stage1_c54_s_fa1;
    wire stage1_c54_c_fa1;
    wire stage1_c54_s_fa2;
    wire stage1_c54_c_fa2;
    wire stage1_c54_s_fa3;
    wire stage1_c54_c_fa3;
    wire stage1_c54_s_fa4;
    wire stage1_c54_c_fa4;
    wire stage1_c54_s_fa5;
    wire stage1_c54_c_fa5;
    wire stage1_c54_s_fa6;
    wire stage1_c54_c_fa6;
    wire stage1_c54_s_fa7;
    wire stage1_c54_c_fa7;
    wire stage1_c54_s_fa8;
    wire stage1_c54_c_fa8;
    wire stage1_c54_s_fa9;
    wire stage1_c54_c_fa9;
    wire stage1_c54_s_fa10;
    wire stage1_c54_c_fa10;
    wire stage1_c54_s_fa11;
    wire stage1_c54_c_fa11;
    wire stage1_c54_s_fa12;
    wire stage1_c54_c_fa12;
    wire stage1_c54_s_ha0;
    wire stage1_c54_c_ha0;
    wire stage1_c55_s_fa0;
    wire stage1_c55_c_fa0;
    wire stage1_c55_s_fa1;
    wire stage1_c55_c_fa1;
    wire stage1_c55_s_fa2;
    wire stage1_c55_c_fa2;
    wire stage1_c55_s_fa3;
    wire stage1_c55_c_fa3;
    wire stage1_c55_s_fa4;
    wire stage1_c55_c_fa4;
    wire stage1_c55_s_fa5;
    wire stage1_c55_c_fa5;
    wire stage1_c55_s_fa6;
    wire stage1_c55_c_fa6;
    wire stage1_c55_s_fa7;
    wire stage1_c55_c_fa7;
    wire stage1_c55_s_fa8;
    wire stage1_c55_c_fa8;
    wire stage1_c55_s_fa9;
    wire stage1_c55_c_fa9;
    wire stage1_c55_s_fa10;
    wire stage1_c55_c_fa10;
    wire stage1_c55_s_fa11;
    wire stage1_c55_c_fa11;
    wire stage1_c55_s_fa12;
    wire stage1_c55_c_fa12;
    wire stage1_c55_s_ha0;
    wire stage1_c55_c_ha0;
    wire stage1_c56_s_fa0;
    wire stage1_c56_c_fa0;
    wire stage1_c56_s_fa1;
    wire stage1_c56_c_fa1;
    wire stage1_c56_s_fa2;
    wire stage1_c56_c_fa2;
    wire stage1_c56_s_fa3;
    wire stage1_c56_c_fa3;
    wire stage1_c56_s_fa4;
    wire stage1_c56_c_fa4;
    wire stage1_c56_s_fa5;
    wire stage1_c56_c_fa5;
    wire stage1_c56_s_fa6;
    wire stage1_c56_c_fa6;
    wire stage1_c56_s_fa7;
    wire stage1_c56_c_fa7;
    wire stage1_c56_s_fa8;
    wire stage1_c56_c_fa8;
    wire stage1_c56_s_fa9;
    wire stage1_c56_c_fa9;
    wire stage1_c56_s_fa10;
    wire stage1_c56_c_fa10;
    wire stage1_c56_s_fa11;
    wire stage1_c56_c_fa11;
    wire stage1_c56_s_fa12;
    wire stage1_c56_c_fa12;
    wire stage1_c56_s_ha0;
    wire stage1_c56_c_ha0;
    wire stage1_c57_s_fa0;
    wire stage1_c57_c_fa0;
    wire stage1_c57_s_fa1;
    wire stage1_c57_c_fa1;
    wire stage1_c57_s_fa2;
    wire stage1_c57_c_fa2;
    wire stage1_c57_s_fa3;
    wire stage1_c57_c_fa3;
    wire stage1_c57_s_fa4;
    wire stage1_c57_c_fa4;
    wire stage1_c57_s_fa5;
    wire stage1_c57_c_fa5;
    wire stage1_c57_s_fa6;
    wire stage1_c57_c_fa6;
    wire stage1_c57_s_fa7;
    wire stage1_c57_c_fa7;
    wire stage1_c57_s_fa8;
    wire stage1_c57_c_fa8;
    wire stage1_c57_s_fa9;
    wire stage1_c57_c_fa9;
    wire stage1_c57_s_fa10;
    wire stage1_c57_c_fa10;
    wire stage1_c57_s_fa11;
    wire stage1_c57_c_fa11;
    wire stage1_c57_s_fa12;
    wire stage1_c57_c_fa12;
    wire stage1_c57_s_ha0;
    wire stage1_c57_c_ha0;
    wire stage1_c58_s_fa0;
    wire stage1_c58_c_fa0;
    wire stage1_c58_s_fa1;
    wire stage1_c58_c_fa1;
    wire stage1_c58_s_fa2;
    wire stage1_c58_c_fa2;
    wire stage1_c58_s_fa3;
    wire stage1_c58_c_fa3;
    wire stage1_c58_s_fa4;
    wire stage1_c58_c_fa4;
    wire stage1_c58_s_fa5;
    wire stage1_c58_c_fa5;
    wire stage1_c58_s_fa6;
    wire stage1_c58_c_fa6;
    wire stage1_c58_s_fa7;
    wire stage1_c58_c_fa7;
    wire stage1_c58_s_fa8;
    wire stage1_c58_c_fa8;
    wire stage1_c58_s_fa9;
    wire stage1_c58_c_fa9;
    wire stage1_c58_s_fa10;
    wire stage1_c58_c_fa10;
    wire stage1_c58_s_fa11;
    wire stage1_c58_c_fa11;
    wire stage1_c58_s_fa12;
    wire stage1_c58_c_fa12;
    wire stage1_c58_s_ha0;
    wire stage1_c58_c_ha0;
    wire stage1_c59_s_fa0;
    wire stage1_c59_c_fa0;
    wire stage1_c59_s_fa1;
    wire stage1_c59_c_fa1;
    wire stage1_c59_s_fa2;
    wire stage1_c59_c_fa2;
    wire stage1_c59_s_fa3;
    wire stage1_c59_c_fa3;
    wire stage1_c59_s_fa4;
    wire stage1_c59_c_fa4;
    wire stage1_c59_s_fa5;
    wire stage1_c59_c_fa5;
    wire stage1_c59_s_fa6;
    wire stage1_c59_c_fa6;
    wire stage1_c59_s_fa7;
    wire stage1_c59_c_fa7;
    wire stage1_c59_s_fa8;
    wire stage1_c59_c_fa8;
    wire stage1_c59_s_fa9;
    wire stage1_c59_c_fa9;
    wire stage1_c59_s_fa10;
    wire stage1_c59_c_fa10;
    wire stage1_c59_s_fa11;
    wire stage1_c59_c_fa11;
    wire stage1_c59_s_fa12;
    wire stage1_c59_c_fa12;
    wire stage1_c59_s_ha0;
    wire stage1_c59_c_ha0;
    wire stage1_c60_s_fa0;
    wire stage1_c60_c_fa0;
    wire stage1_c60_s_fa1;
    wire stage1_c60_c_fa1;
    wire stage1_c60_s_fa2;
    wire stage1_c60_c_fa2;
    wire stage1_c60_s_fa3;
    wire stage1_c60_c_fa3;
    wire stage1_c60_s_fa4;
    wire stage1_c60_c_fa4;
    wire stage1_c60_s_fa5;
    wire stage1_c60_c_fa5;
    wire stage1_c60_s_fa6;
    wire stage1_c60_c_fa6;
    wire stage1_c60_s_fa7;
    wire stage1_c60_c_fa7;
    wire stage1_c60_s_fa8;
    wire stage1_c60_c_fa8;
    wire stage1_c60_s_fa9;
    wire stage1_c60_c_fa9;
    wire stage1_c60_s_fa10;
    wire stage1_c60_c_fa10;
    wire stage1_c60_s_fa11;
    wire stage1_c60_c_fa11;
    wire stage1_c60_s_fa12;
    wire stage1_c60_c_fa12;
    wire stage1_c60_s_ha0;
    wire stage1_c60_c_ha0;
    wire stage1_c61_s_fa0;
    wire stage1_c61_c_fa0;
    wire stage1_c61_s_fa1;
    wire stage1_c61_c_fa1;
    wire stage1_c61_s_fa2;
    wire stage1_c61_c_fa2;
    wire stage1_c61_s_fa3;
    wire stage1_c61_c_fa3;
    wire stage1_c61_s_fa4;
    wire stage1_c61_c_fa4;
    wire stage1_c61_s_fa5;
    wire stage1_c61_c_fa5;
    wire stage1_c61_s_fa6;
    wire stage1_c61_c_fa6;
    wire stage1_c61_s_fa7;
    wire stage1_c61_c_fa7;
    wire stage1_c61_s_fa8;
    wire stage1_c61_c_fa8;
    wire stage1_c61_s_fa9;
    wire stage1_c61_c_fa9;
    wire stage1_c61_s_fa10;
    wire stage1_c61_c_fa10;
    wire stage1_c61_s_fa11;
    wire stage1_c61_c_fa11;
    wire stage1_c61_s_fa12;
    wire stage1_c61_c_fa12;
    wire stage1_c61_s_ha0;
    wire stage1_c61_c_ha0;
    wire stage1_c62_s_fa0;
    wire stage1_c62_c_fa0;
    wire stage1_c62_s_fa1;
    wire stage1_c62_c_fa1;
    wire stage1_c62_s_fa2;
    wire stage1_c62_c_fa2;
    wire stage1_c62_s_fa3;
    wire stage1_c62_c_fa3;
    wire stage1_c62_s_fa4;
    wire stage1_c62_c_fa4;
    wire stage1_c62_s_fa5;
    wire stage1_c62_c_fa5;
    wire stage1_c62_s_fa6;
    wire stage1_c62_c_fa6;
    wire stage1_c62_s_fa7;
    wire stage1_c62_c_fa7;
    wire stage1_c62_s_fa8;
    wire stage1_c62_c_fa8;
    wire stage1_c62_s_fa9;
    wire stage1_c62_c_fa9;
    wire stage1_c62_s_fa10;
    wire stage1_c62_c_fa10;
    wire stage1_c62_s_fa11;
    wire stage1_c62_c_fa11;
    wire stage1_c62_s_fa12;
    wire stage1_c62_c_fa12;
    wire stage1_c62_s_ha0;
    wire stage1_c62_c_ha0;
    wire stage1_c63_s_fa0;
    wire stage1_c63_c_fa0;
    wire stage1_c63_s_fa1;
    wire stage1_c63_c_fa1;
    wire stage1_c63_s_fa2;
    wire stage1_c63_c_fa2;
    wire stage1_c63_s_fa3;
    wire stage1_c63_c_fa3;
    wire stage1_c63_s_fa4;
    wire stage1_c63_c_fa4;
    wire stage1_c63_s_fa5;
    wire stage1_c63_c_fa5;
    wire stage1_c63_s_fa6;
    wire stage1_c63_c_fa6;
    wire stage1_c63_s_fa7;
    wire stage1_c63_c_fa7;
    wire stage1_c63_s_fa8;
    wire stage1_c63_c_fa8;
    wire stage1_c63_s_fa9;
    wire stage1_c63_c_fa9;
    wire stage1_c63_s_fa10;
    wire stage1_c63_c_fa10;
    wire stage1_c63_s_fa11;
    wire stage1_c63_c_fa11;
    wire stage1_c63_s_fa12;
    wire stage1_c63_c_fa12;
    wire stage1_c63_s_ha0;
    wire stage1_c63_c_ha0;
    wire stage1_c64_s_fa0;
    wire stage1_c64_c_fa0;
    wire stage1_c64_s_fa1;
    wire stage1_c64_c_fa1;
    wire stage1_c64_s_fa2;
    wire stage1_c64_c_fa2;
    wire stage1_c64_s_fa3;
    wire stage1_c64_c_fa3;
    wire stage1_c64_s_fa4;
    wire stage1_c64_c_fa4;
    wire stage1_c64_s_fa5;
    wire stage1_c64_c_fa5;
    wire stage1_c64_s_fa6;
    wire stage1_c64_c_fa6;
    wire stage1_c64_s_fa7;
    wire stage1_c64_c_fa7;
    wire stage1_c64_s_fa8;
    wire stage1_c64_c_fa8;
    wire stage1_c64_s_fa9;
    wire stage1_c64_c_fa9;
    wire stage1_c64_s_fa10;
    wire stage1_c64_c_fa10;
    wire stage1_c64_s_fa11;
    wire stage1_c64_c_fa11;
    wire stage1_c64_s_fa12;
    wire stage1_c64_c_fa12;
    wire stage1_c64_s_ha0;
    wire stage1_c64_c_ha0;
    wire stage1_c65_s_fa0;
    wire stage1_c65_c_fa0;
    wire stage1_c65_s_fa1;
    wire stage1_c65_c_fa1;
    wire stage1_c65_s_fa2;
    wire stage1_c65_c_fa2;
    wire stage1_c65_s_fa3;
    wire stage1_c65_c_fa3;
    wire stage1_c65_s_fa4;
    wire stage1_c65_c_fa4;
    wire stage1_c65_s_fa5;
    wire stage1_c65_c_fa5;
    wire stage1_c65_s_fa6;
    wire stage1_c65_c_fa6;
    wire stage1_c65_s_fa7;
    wire stage1_c65_c_fa7;
    wire stage1_c65_s_fa8;
    wire stage1_c65_c_fa8;
    wire stage1_c65_s_fa9;
    wire stage1_c65_c_fa9;
    wire stage1_c65_s_fa10;
    wire stage1_c65_c_fa10;
    wire stage1_c65_s_fa11;
    wire stage1_c65_c_fa11;
    wire stage1_c65_s_fa12;
    wire stage1_c65_c_fa12;
    wire stage1_c65_s_ha0;
    wire stage1_c65_c_ha0;
    wire stage1_c66_s_fa0;
    wire stage1_c66_c_fa0;
    wire stage1_c66_s_fa1;
    wire stage1_c66_c_fa1;
    wire stage1_c66_s_fa2;
    wire stage1_c66_c_fa2;
    wire stage1_c66_s_fa3;
    wire stage1_c66_c_fa3;
    wire stage1_c66_s_fa4;
    wire stage1_c66_c_fa4;
    wire stage1_c66_s_fa5;
    wire stage1_c66_c_fa5;
    wire stage1_c66_s_fa6;
    wire stage1_c66_c_fa6;
    wire stage1_c66_s_fa7;
    wire stage1_c66_c_fa7;
    wire stage1_c66_s_fa8;
    wire stage1_c66_c_fa8;
    wire stage1_c66_s_fa9;
    wire stage1_c66_c_fa9;
    wire stage1_c66_s_fa10;
    wire stage1_c66_c_fa10;
    wire stage1_c66_s_fa11;
    wire stage1_c66_c_fa11;
    wire stage1_c66_s_fa12;
    wire stage1_c66_c_fa12;
    wire stage1_c66_s_ha0;
    wire stage1_c66_c_ha0;
    wire stage1_c67_s_fa0;
    wire stage1_c67_c_fa0;
    wire stage1_c67_s_fa1;
    wire stage1_c67_c_fa1;
    wire stage1_c67_s_fa2;
    wire stage1_c67_c_fa2;
    wire stage1_c67_s_fa3;
    wire stage1_c67_c_fa3;
    wire stage1_c67_s_fa4;
    wire stage1_c67_c_fa4;
    wire stage1_c67_s_fa5;
    wire stage1_c67_c_fa5;
    wire stage1_c67_s_fa6;
    wire stage1_c67_c_fa6;
    wire stage1_c67_s_fa7;
    wire stage1_c67_c_fa7;
    wire stage1_c67_s_fa8;
    wire stage1_c67_c_fa8;
    wire stage1_c67_s_fa9;
    wire stage1_c67_c_fa9;
    wire stage1_c67_s_fa10;
    wire stage1_c67_c_fa10;
    wire stage1_c67_s_fa11;
    wire stage1_c67_c_fa11;
    wire stage1_c67_s_fa12;
    wire stage1_c67_c_fa12;
    wire stage1_c67_s_ha0;
    wire stage1_c67_c_ha0;
    wire stage1_c68_s_fa0;
    wire stage1_c68_c_fa0;
    wire stage1_c68_s_fa1;
    wire stage1_c68_c_fa1;
    wire stage1_c68_s_fa2;
    wire stage1_c68_c_fa2;
    wire stage1_c68_s_fa3;
    wire stage1_c68_c_fa3;
    wire stage1_c68_s_fa4;
    wire stage1_c68_c_fa4;
    wire stage1_c68_s_fa5;
    wire stage1_c68_c_fa5;
    wire stage1_c68_s_fa6;
    wire stage1_c68_c_fa6;
    wire stage1_c68_s_fa7;
    wire stage1_c68_c_fa7;
    wire stage1_c68_s_fa8;
    wire stage1_c68_c_fa8;
    wire stage1_c68_s_fa9;
    wire stage1_c68_c_fa9;
    wire stage1_c68_s_fa10;
    wire stage1_c68_c_fa10;
    wire stage1_c68_s_fa11;
    wire stage1_c68_c_fa11;
    wire stage1_c68_s_fa12;
    wire stage1_c68_c_fa12;
    wire stage1_c68_s_ha0;
    wire stage1_c68_c_ha0;
    wire stage1_c69_s_fa0;
    wire stage1_c69_c_fa0;
    wire stage1_c69_s_fa1;
    wire stage1_c69_c_fa1;
    wire stage1_c69_s_fa2;
    wire stage1_c69_c_fa2;
    wire stage1_c69_s_fa3;
    wire stage1_c69_c_fa3;
    wire stage1_c69_s_fa4;
    wire stage1_c69_c_fa4;
    wire stage1_c69_s_fa5;
    wire stage1_c69_c_fa5;
    wire stage1_c69_s_fa6;
    wire stage1_c69_c_fa6;
    wire stage1_c69_s_fa7;
    wire stage1_c69_c_fa7;
    wire stage1_c69_s_fa8;
    wire stage1_c69_c_fa8;
    wire stage1_c69_s_fa9;
    wire stage1_c69_c_fa9;
    wire stage1_c69_s_fa10;
    wire stage1_c69_c_fa10;
    wire stage1_c69_s_fa11;
    wire stage1_c69_c_fa11;
    wire stage1_c69_s_fa12;
    wire stage1_c69_c_fa12;
    wire stage1_c69_s_ha0;
    wire stage1_c69_c_ha0;
    wire stage1_c70_s_fa0;
    wire stage1_c70_c_fa0;
    wire stage1_c70_s_fa1;
    wire stage1_c70_c_fa1;
    wire stage1_c70_s_fa2;
    wire stage1_c70_c_fa2;
    wire stage1_c70_s_fa3;
    wire stage1_c70_c_fa3;
    wire stage1_c70_s_fa4;
    wire stage1_c70_c_fa4;
    wire stage1_c70_s_fa5;
    wire stage1_c70_c_fa5;
    wire stage1_c70_s_fa6;
    wire stage1_c70_c_fa6;
    wire stage1_c70_s_fa7;
    wire stage1_c70_c_fa7;
    wire stage1_c70_s_fa8;
    wire stage1_c70_c_fa8;
    wire stage1_c70_s_fa9;
    wire stage1_c70_c_fa9;
    wire stage1_c70_s_fa10;
    wire stage1_c70_c_fa10;
    wire stage1_c70_s_fa11;
    wire stage1_c70_c_fa11;
    wire stage1_c70_s_fa12;
    wire stage1_c70_c_fa12;
    wire stage1_c70_s_ha0;
    wire stage1_c70_c_ha0;
    wire stage1_c71_s_fa0;
    wire stage1_c71_c_fa0;
    wire stage1_c71_s_fa1;
    wire stage1_c71_c_fa1;
    wire stage1_c71_s_fa2;
    wire stage1_c71_c_fa2;
    wire stage1_c71_s_fa3;
    wire stage1_c71_c_fa3;
    wire stage1_c71_s_fa4;
    wire stage1_c71_c_fa4;
    wire stage1_c71_s_fa5;
    wire stage1_c71_c_fa5;
    wire stage1_c71_s_fa6;
    wire stage1_c71_c_fa6;
    wire stage1_c71_s_fa7;
    wire stage1_c71_c_fa7;
    wire stage1_c71_s_fa8;
    wire stage1_c71_c_fa8;
    wire stage1_c71_s_fa9;
    wire stage1_c71_c_fa9;
    wire stage1_c71_s_fa10;
    wire stage1_c71_c_fa10;
    wire stage1_c71_s_fa11;
    wire stage1_c71_c_fa11;
    wire stage1_c71_s_fa12;
    wire stage1_c71_c_fa12;
    wire stage1_c71_s_ha0;
    wire stage1_c71_c_ha0;
    wire stage1_c72_s_fa0;
    wire stage1_c72_c_fa0;
    wire stage1_c72_s_fa1;
    wire stage1_c72_c_fa1;
    wire stage1_c72_s_fa2;
    wire stage1_c72_c_fa2;
    wire stage1_c72_s_fa3;
    wire stage1_c72_c_fa3;
    wire stage1_c72_s_fa4;
    wire stage1_c72_c_fa4;
    wire stage1_c72_s_fa5;
    wire stage1_c72_c_fa5;
    wire stage1_c72_s_fa6;
    wire stage1_c72_c_fa6;
    wire stage1_c72_s_fa7;
    wire stage1_c72_c_fa7;
    wire stage1_c72_s_fa8;
    wire stage1_c72_c_fa8;
    wire stage1_c72_s_fa9;
    wire stage1_c72_c_fa9;
    wire stage1_c72_s_fa10;
    wire stage1_c72_c_fa10;
    wire stage1_c72_s_fa11;
    wire stage1_c72_c_fa11;
    wire stage1_c72_s_fa12;
    wire stage1_c72_c_fa12;
    wire stage1_c73_s_fa0;
    wire stage1_c73_c_fa0;
    wire stage1_c73_s_fa1;
    wire stage1_c73_c_fa1;
    wire stage1_c73_s_fa2;
    wire stage1_c73_c_fa2;
    wire stage1_c73_s_fa3;
    wire stage1_c73_c_fa3;
    wire stage1_c73_s_fa4;
    wire stage1_c73_c_fa4;
    wire stage1_c73_s_fa5;
    wire stage1_c73_c_fa5;
    wire stage1_c73_s_fa6;
    wire stage1_c73_c_fa6;
    wire stage1_c73_s_fa7;
    wire stage1_c73_c_fa7;
    wire stage1_c73_s_fa8;
    wire stage1_c73_c_fa8;
    wire stage1_c73_s_fa9;
    wire stage1_c73_c_fa9;
    wire stage1_c73_s_fa10;
    wire stage1_c73_c_fa10;
    wire stage1_c73_s_fa11;
    wire stage1_c73_c_fa11;
    wire stage1_c73_s_fa12;
    wire stage1_c73_c_fa12;
    wire stage1_c74_s_fa0;
    wire stage1_c74_c_fa0;
    wire stage1_c74_s_fa1;
    wire stage1_c74_c_fa1;
    wire stage1_c74_s_fa2;
    wire stage1_c74_c_fa2;
    wire stage1_c74_s_fa3;
    wire stage1_c74_c_fa3;
    wire stage1_c74_s_fa4;
    wire stage1_c74_c_fa4;
    wire stage1_c74_s_fa5;
    wire stage1_c74_c_fa5;
    wire stage1_c74_s_fa6;
    wire stage1_c74_c_fa6;
    wire stage1_c74_s_fa7;
    wire stage1_c74_c_fa7;
    wire stage1_c74_s_fa8;
    wire stage1_c74_c_fa8;
    wire stage1_c74_s_fa9;
    wire stage1_c74_c_fa9;
    wire stage1_c74_s_fa10;
    wire stage1_c74_c_fa10;
    wire stage1_c74_s_fa11;
    wire stage1_c74_c_fa11;
    wire stage1_c74_s_ha0;
    wire stage1_c74_c_ha0;
    wire stage1_c75_s_fa0;
    wire stage1_c75_c_fa0;
    wire stage1_c75_s_fa1;
    wire stage1_c75_c_fa1;
    wire stage1_c75_s_fa2;
    wire stage1_c75_c_fa2;
    wire stage1_c75_s_fa3;
    wire stage1_c75_c_fa3;
    wire stage1_c75_s_fa4;
    wire stage1_c75_c_fa4;
    wire stage1_c75_s_fa5;
    wire stage1_c75_c_fa5;
    wire stage1_c75_s_fa6;
    wire stage1_c75_c_fa6;
    wire stage1_c75_s_fa7;
    wire stage1_c75_c_fa7;
    wire stage1_c75_s_fa8;
    wire stage1_c75_c_fa8;
    wire stage1_c75_s_fa9;
    wire stage1_c75_c_fa9;
    wire stage1_c75_s_fa10;
    wire stage1_c75_c_fa10;
    wire stage1_c75_s_fa11;
    wire stage1_c75_c_fa11;
    wire stage1_c76_s_fa0;
    wire stage1_c76_c_fa0;
    wire stage1_c76_s_fa1;
    wire stage1_c76_c_fa1;
    wire stage1_c76_s_fa2;
    wire stage1_c76_c_fa2;
    wire stage1_c76_s_fa3;
    wire stage1_c76_c_fa3;
    wire stage1_c76_s_fa4;
    wire stage1_c76_c_fa4;
    wire stage1_c76_s_fa5;
    wire stage1_c76_c_fa5;
    wire stage1_c76_s_fa6;
    wire stage1_c76_c_fa6;
    wire stage1_c76_s_fa7;
    wire stage1_c76_c_fa7;
    wire stage1_c76_s_fa8;
    wire stage1_c76_c_fa8;
    wire stage1_c76_s_fa9;
    wire stage1_c76_c_fa9;
    wire stage1_c76_s_fa10;
    wire stage1_c76_c_fa10;
    wire stage1_c76_s_fa11;
    wire stage1_c76_c_fa11;
    wire stage1_c77_s_fa0;
    wire stage1_c77_c_fa0;
    wire stage1_c77_s_fa1;
    wire stage1_c77_c_fa1;
    wire stage1_c77_s_fa2;
    wire stage1_c77_c_fa2;
    wire stage1_c77_s_fa3;
    wire stage1_c77_c_fa3;
    wire stage1_c77_s_fa4;
    wire stage1_c77_c_fa4;
    wire stage1_c77_s_fa5;
    wire stage1_c77_c_fa5;
    wire stage1_c77_s_fa6;
    wire stage1_c77_c_fa6;
    wire stage1_c77_s_fa7;
    wire stage1_c77_c_fa7;
    wire stage1_c77_s_fa8;
    wire stage1_c77_c_fa8;
    wire stage1_c77_s_fa9;
    wire stage1_c77_c_fa9;
    wire stage1_c77_s_fa10;
    wire stage1_c77_c_fa10;
    wire stage1_c77_s_ha0;
    wire stage1_c77_c_ha0;
    wire stage1_c78_s_fa0;
    wire stage1_c78_c_fa0;
    wire stage1_c78_s_fa1;
    wire stage1_c78_c_fa1;
    wire stage1_c78_s_fa2;
    wire stage1_c78_c_fa2;
    wire stage1_c78_s_fa3;
    wire stage1_c78_c_fa3;
    wire stage1_c78_s_fa4;
    wire stage1_c78_c_fa4;
    wire stage1_c78_s_fa5;
    wire stage1_c78_c_fa5;
    wire stage1_c78_s_fa6;
    wire stage1_c78_c_fa6;
    wire stage1_c78_s_fa7;
    wire stage1_c78_c_fa7;
    wire stage1_c78_s_fa8;
    wire stage1_c78_c_fa8;
    wire stage1_c78_s_fa9;
    wire stage1_c78_c_fa9;
    wire stage1_c78_s_fa10;
    wire stage1_c78_c_fa10;
    wire stage1_c79_s_fa0;
    wire stage1_c79_c_fa0;
    wire stage1_c79_s_fa1;
    wire stage1_c79_c_fa1;
    wire stage1_c79_s_fa2;
    wire stage1_c79_c_fa2;
    wire stage1_c79_s_fa3;
    wire stage1_c79_c_fa3;
    wire stage1_c79_s_fa4;
    wire stage1_c79_c_fa4;
    wire stage1_c79_s_fa5;
    wire stage1_c79_c_fa5;
    wire stage1_c79_s_fa6;
    wire stage1_c79_c_fa6;
    wire stage1_c79_s_fa7;
    wire stage1_c79_c_fa7;
    wire stage1_c79_s_fa8;
    wire stage1_c79_c_fa8;
    wire stage1_c79_s_fa9;
    wire stage1_c79_c_fa9;
    wire stage1_c79_s_fa10;
    wire stage1_c79_c_fa10;
    wire stage1_c80_s_fa0;
    wire stage1_c80_c_fa0;
    wire stage1_c80_s_fa1;
    wire stage1_c80_c_fa1;
    wire stage1_c80_s_fa2;
    wire stage1_c80_c_fa2;
    wire stage1_c80_s_fa3;
    wire stage1_c80_c_fa3;
    wire stage1_c80_s_fa4;
    wire stage1_c80_c_fa4;
    wire stage1_c80_s_fa5;
    wire stage1_c80_c_fa5;
    wire stage1_c80_s_fa6;
    wire stage1_c80_c_fa6;
    wire stage1_c80_s_fa7;
    wire stage1_c80_c_fa7;
    wire stage1_c80_s_fa8;
    wire stage1_c80_c_fa8;
    wire stage1_c80_s_fa9;
    wire stage1_c80_c_fa9;
    wire stage1_c80_s_ha0;
    wire stage1_c80_c_ha0;
    wire stage1_c81_s_fa0;
    wire stage1_c81_c_fa0;
    wire stage1_c81_s_fa1;
    wire stage1_c81_c_fa1;
    wire stage1_c81_s_fa2;
    wire stage1_c81_c_fa2;
    wire stage1_c81_s_fa3;
    wire stage1_c81_c_fa3;
    wire stage1_c81_s_fa4;
    wire stage1_c81_c_fa4;
    wire stage1_c81_s_fa5;
    wire stage1_c81_c_fa5;
    wire stage1_c81_s_fa6;
    wire stage1_c81_c_fa6;
    wire stage1_c81_s_fa7;
    wire stage1_c81_c_fa7;
    wire stage1_c81_s_fa8;
    wire stage1_c81_c_fa8;
    wire stage1_c81_s_fa9;
    wire stage1_c81_c_fa9;
    wire stage1_c82_s_fa0;
    wire stage1_c82_c_fa0;
    wire stage1_c82_s_fa1;
    wire stage1_c82_c_fa1;
    wire stage1_c82_s_fa2;
    wire stage1_c82_c_fa2;
    wire stage1_c82_s_fa3;
    wire stage1_c82_c_fa3;
    wire stage1_c82_s_fa4;
    wire stage1_c82_c_fa4;
    wire stage1_c82_s_fa5;
    wire stage1_c82_c_fa5;
    wire stage1_c82_s_fa6;
    wire stage1_c82_c_fa6;
    wire stage1_c82_s_fa7;
    wire stage1_c82_c_fa7;
    wire stage1_c82_s_fa8;
    wire stage1_c82_c_fa8;
    wire stage1_c82_s_fa9;
    wire stage1_c82_c_fa9;
    wire stage1_c83_s_fa0;
    wire stage1_c83_c_fa0;
    wire stage1_c83_s_fa1;
    wire stage1_c83_c_fa1;
    wire stage1_c83_s_fa2;
    wire stage1_c83_c_fa2;
    wire stage1_c83_s_fa3;
    wire stage1_c83_c_fa3;
    wire stage1_c83_s_fa4;
    wire stage1_c83_c_fa4;
    wire stage1_c83_s_fa5;
    wire stage1_c83_c_fa5;
    wire stage1_c83_s_fa6;
    wire stage1_c83_c_fa6;
    wire stage1_c83_s_fa7;
    wire stage1_c83_c_fa7;
    wire stage1_c83_s_fa8;
    wire stage1_c83_c_fa8;
    wire stage1_c83_s_ha0;
    wire stage1_c83_c_ha0;
    wire stage1_c84_s_fa0;
    wire stage1_c84_c_fa0;
    wire stage1_c84_s_fa1;
    wire stage1_c84_c_fa1;
    wire stage1_c84_s_fa2;
    wire stage1_c84_c_fa2;
    wire stage1_c84_s_fa3;
    wire stage1_c84_c_fa3;
    wire stage1_c84_s_fa4;
    wire stage1_c84_c_fa4;
    wire stage1_c84_s_fa5;
    wire stage1_c84_c_fa5;
    wire stage1_c84_s_fa6;
    wire stage1_c84_c_fa6;
    wire stage1_c84_s_fa7;
    wire stage1_c84_c_fa7;
    wire stage1_c84_s_fa8;
    wire stage1_c84_c_fa8;
    wire stage1_c85_s_fa0;
    wire stage1_c85_c_fa0;
    wire stage1_c85_s_fa1;
    wire stage1_c85_c_fa1;
    wire stage1_c85_s_fa2;
    wire stage1_c85_c_fa2;
    wire stage1_c85_s_fa3;
    wire stage1_c85_c_fa3;
    wire stage1_c85_s_fa4;
    wire stage1_c85_c_fa4;
    wire stage1_c85_s_fa5;
    wire stage1_c85_c_fa5;
    wire stage1_c85_s_fa6;
    wire stage1_c85_c_fa6;
    wire stage1_c85_s_fa7;
    wire stage1_c85_c_fa7;
    wire stage1_c85_s_fa8;
    wire stage1_c85_c_fa8;
    wire stage1_c86_s_fa0;
    wire stage1_c86_c_fa0;
    wire stage1_c86_s_fa1;
    wire stage1_c86_c_fa1;
    wire stage1_c86_s_fa2;
    wire stage1_c86_c_fa2;
    wire stage1_c86_s_fa3;
    wire stage1_c86_c_fa3;
    wire stage1_c86_s_fa4;
    wire stage1_c86_c_fa4;
    wire stage1_c86_s_fa5;
    wire stage1_c86_c_fa5;
    wire stage1_c86_s_fa6;
    wire stage1_c86_c_fa6;
    wire stage1_c86_s_fa7;
    wire stage1_c86_c_fa7;
    wire stage1_c86_s_ha0;
    wire stage1_c86_c_ha0;
    wire stage1_c87_s_fa0;
    wire stage1_c87_c_fa0;
    wire stage1_c87_s_fa1;
    wire stage1_c87_c_fa1;
    wire stage1_c87_s_fa2;
    wire stage1_c87_c_fa2;
    wire stage1_c87_s_fa3;
    wire stage1_c87_c_fa3;
    wire stage1_c87_s_fa4;
    wire stage1_c87_c_fa4;
    wire stage1_c87_s_fa5;
    wire stage1_c87_c_fa5;
    wire stage1_c87_s_fa6;
    wire stage1_c87_c_fa6;
    wire stage1_c87_s_fa7;
    wire stage1_c87_c_fa7;
    wire stage1_c88_s_fa0;
    wire stage1_c88_c_fa0;
    wire stage1_c88_s_fa1;
    wire stage1_c88_c_fa1;
    wire stage1_c88_s_fa2;
    wire stage1_c88_c_fa2;
    wire stage1_c88_s_fa3;
    wire stage1_c88_c_fa3;
    wire stage1_c88_s_fa4;
    wire stage1_c88_c_fa4;
    wire stage1_c88_s_fa5;
    wire stage1_c88_c_fa5;
    wire stage1_c88_s_fa6;
    wire stage1_c88_c_fa6;
    wire stage1_c88_s_fa7;
    wire stage1_c88_c_fa7;
    wire stage1_c89_s_fa0;
    wire stage1_c89_c_fa0;
    wire stage1_c89_s_fa1;
    wire stage1_c89_c_fa1;
    wire stage1_c89_s_fa2;
    wire stage1_c89_c_fa2;
    wire stage1_c89_s_fa3;
    wire stage1_c89_c_fa3;
    wire stage1_c89_s_fa4;
    wire stage1_c89_c_fa4;
    wire stage1_c89_s_fa5;
    wire stage1_c89_c_fa5;
    wire stage1_c89_s_fa6;
    wire stage1_c89_c_fa6;
    wire stage1_c89_s_ha0;
    wire stage1_c89_c_ha0;
    wire stage1_c90_s_fa0;
    wire stage1_c90_c_fa0;
    wire stage1_c90_s_fa1;
    wire stage1_c90_c_fa1;
    wire stage1_c90_s_fa2;
    wire stage1_c90_c_fa2;
    wire stage1_c90_s_fa3;
    wire stage1_c90_c_fa3;
    wire stage1_c90_s_fa4;
    wire stage1_c90_c_fa4;
    wire stage1_c90_s_fa5;
    wire stage1_c90_c_fa5;
    wire stage1_c90_s_fa6;
    wire stage1_c90_c_fa6;
    wire stage1_c91_s_fa0;
    wire stage1_c91_c_fa0;
    wire stage1_c91_s_fa1;
    wire stage1_c91_c_fa1;
    wire stage1_c91_s_fa2;
    wire stage1_c91_c_fa2;
    wire stage1_c91_s_fa3;
    wire stage1_c91_c_fa3;
    wire stage1_c91_s_fa4;
    wire stage1_c91_c_fa4;
    wire stage1_c91_s_fa5;
    wire stage1_c91_c_fa5;
    wire stage1_c91_s_fa6;
    wire stage1_c91_c_fa6;
    wire stage1_c92_s_fa0;
    wire stage1_c92_c_fa0;
    wire stage1_c92_s_fa1;
    wire stage1_c92_c_fa1;
    wire stage1_c92_s_fa2;
    wire stage1_c92_c_fa2;
    wire stage1_c92_s_fa3;
    wire stage1_c92_c_fa3;
    wire stage1_c92_s_fa4;
    wire stage1_c92_c_fa4;
    wire stage1_c92_s_fa5;
    wire stage1_c92_c_fa5;
    wire stage1_c92_s_ha0;
    wire stage1_c92_c_ha0;
    wire stage1_c93_s_fa0;
    wire stage1_c93_c_fa0;
    wire stage1_c93_s_fa1;
    wire stage1_c93_c_fa1;
    wire stage1_c93_s_fa2;
    wire stage1_c93_c_fa2;
    wire stage1_c93_s_fa3;
    wire stage1_c93_c_fa3;
    wire stage1_c93_s_fa4;
    wire stage1_c93_c_fa4;
    wire stage1_c93_s_fa5;
    wire stage1_c93_c_fa5;
    wire stage1_c94_s_fa0;
    wire stage1_c94_c_fa0;
    wire stage1_c94_s_fa1;
    wire stage1_c94_c_fa1;
    wire stage1_c94_s_fa2;
    wire stage1_c94_c_fa2;
    wire stage1_c94_s_fa3;
    wire stage1_c94_c_fa3;
    wire stage1_c94_s_fa4;
    wire stage1_c94_c_fa4;
    wire stage1_c94_s_fa5;
    wire stage1_c94_c_fa5;
    wire stage1_c95_s_fa0;
    wire stage1_c95_c_fa0;
    wire stage1_c95_s_fa1;
    wire stage1_c95_c_fa1;
    wire stage1_c95_s_fa2;
    wire stage1_c95_c_fa2;
    wire stage1_c95_s_fa3;
    wire stage1_c95_c_fa3;
    wire stage1_c95_s_fa4;
    wire stage1_c95_c_fa4;
    wire stage1_c95_s_ha0;
    wire stage1_c95_c_ha0;
    wire stage1_c96_s_fa0;
    wire stage1_c96_c_fa0;
    wire stage1_c96_s_fa1;
    wire stage1_c96_c_fa1;
    wire stage1_c96_s_fa2;
    wire stage1_c96_c_fa2;
    wire stage1_c96_s_fa3;
    wire stage1_c96_c_fa3;
    wire stage1_c96_s_fa4;
    wire stage1_c96_c_fa4;
    wire stage1_c97_s_fa0;
    wire stage1_c97_c_fa0;
    wire stage1_c97_s_fa1;
    wire stage1_c97_c_fa1;
    wire stage1_c97_s_fa2;
    wire stage1_c97_c_fa2;
    wire stage1_c97_s_fa3;
    wire stage1_c97_c_fa3;
    wire stage1_c97_s_fa4;
    wire stage1_c97_c_fa4;
    wire stage1_c98_s_fa0;
    wire stage1_c98_c_fa0;
    wire stage1_c98_s_fa1;
    wire stage1_c98_c_fa1;
    wire stage1_c98_s_fa2;
    wire stage1_c98_c_fa2;
    wire stage1_c98_s_fa3;
    wire stage1_c98_c_fa3;
    wire stage1_c98_s_ha0;
    wire stage1_c98_c_ha0;
    wire stage1_c99_s_fa0;
    wire stage1_c99_c_fa0;
    wire stage1_c99_s_fa1;
    wire stage1_c99_c_fa1;
    wire stage1_c99_s_fa2;
    wire stage1_c99_c_fa2;
    wire stage1_c99_s_fa3;
    wire stage1_c99_c_fa3;
    wire stage1_c100_s_fa0;
    wire stage1_c100_c_fa0;
    wire stage1_c100_s_fa1;
    wire stage1_c100_c_fa1;
    wire stage1_c100_s_fa2;
    wire stage1_c100_c_fa2;
    wire stage1_c100_s_fa3;
    wire stage1_c100_c_fa3;
    wire stage1_c101_s_fa0;
    wire stage1_c101_c_fa0;
    wire stage1_c101_s_fa1;
    wire stage1_c101_c_fa1;
    wire stage1_c101_s_fa2;
    wire stage1_c101_c_fa2;
    wire stage1_c101_s_ha0;
    wire stage1_c101_c_ha0;
    wire stage1_c102_s_fa0;
    wire stage1_c102_c_fa0;
    wire stage1_c102_s_fa1;
    wire stage1_c102_c_fa1;
    wire stage1_c102_s_fa2;
    wire stage1_c102_c_fa2;
    wire stage1_c103_s_fa0;
    wire stage1_c103_c_fa0;
    wire stage1_c103_s_fa1;
    wire stage1_c103_c_fa1;
    wire stage1_c103_s_fa2;
    wire stage1_c103_c_fa2;
    wire stage1_c104_s_fa0;
    wire stage1_c104_c_fa0;
    wire stage1_c104_s_fa1;
    wire stage1_c104_c_fa1;
    wire stage1_c104_s_ha0;
    wire stage1_c104_c_ha0;
    wire stage1_c105_s_fa0;
    wire stage1_c105_c_fa0;
    wire stage1_c105_s_fa1;
    wire stage1_c105_c_fa1;
    wire stage1_c106_s_fa0;
    wire stage1_c106_c_fa0;
    wire stage1_c106_s_fa1;
    wire stage1_c106_c_fa1;
    wire stage1_c107_s_fa0;
    wire stage1_c107_c_fa0;
    wire stage1_c107_s_ha0;
    wire stage1_c107_c_ha0;
    wire stage1_c108_s_fa0;
    wire stage1_c108_c_fa0;
    wire stage1_c109_s_fa0;
    wire stage1_c109_c_fa0;
    wire stage1_c110_s_ha0;
    wire stage1_c110_c_ha0;
    wire stage2_c2_s_ha0;
    wire stage2_c2_c_ha0;
    wire stage2_c3_s_fa0;
    wire stage2_c3_c_fa0;
    wire stage2_c4_s_fa0;
    wire stage2_c4_c_fa0;
    wire stage2_c5_s_fa0;
    wire stage2_c5_c_fa0;
    wire stage2_c6_s_fa0;
    wire stage2_c6_c_fa0;
    wire stage2_c6_s_ha0;
    wire stage2_c6_c_ha0;
    wire stage2_c7_s_fa0;
    wire stage2_c7_c_fa0;
    wire stage2_c7_s_ha0;
    wire stage2_c7_c_ha0;
    wire stage2_c8_s_fa0;
    wire stage2_c8_c_fa0;
    wire stage2_c8_s_fa1;
    wire stage2_c8_c_fa1;
    wire stage2_c9_s_fa0;
    wire stage2_c9_c_fa0;
    wire stage2_c9_s_fa1;
    wire stage2_c9_c_fa1;
    wire stage2_c10_s_fa0;
    wire stage2_c10_c_fa0;
    wire stage2_c10_s_fa1;
    wire stage2_c10_c_fa1;
    wire stage2_c11_s_fa0;
    wire stage2_c11_c_fa0;
    wire stage2_c11_s_fa1;
    wire stage2_c11_c_fa1;
    wire stage2_c11_s_ha0;
    wire stage2_c11_c_ha0;
    wire stage2_c12_s_fa0;
    wire stage2_c12_c_fa0;
    wire stage2_c12_s_fa1;
    wire stage2_c12_c_fa1;
    wire stage2_c12_s_fa2;
    wire stage2_c12_c_fa2;
    wire stage2_c13_s_fa0;
    wire stage2_c13_c_fa0;
    wire stage2_c13_s_fa1;
    wire stage2_c13_c_fa1;
    wire stage2_c13_s_fa2;
    wire stage2_c13_c_fa2;
    wire stage2_c14_s_fa0;
    wire stage2_c14_c_fa0;
    wire stage2_c14_s_fa1;
    wire stage2_c14_c_fa1;
    wire stage2_c14_s_fa2;
    wire stage2_c14_c_fa2;
    wire stage2_c15_s_fa0;
    wire stage2_c15_c_fa0;
    wire stage2_c15_s_fa1;
    wire stage2_c15_c_fa1;
    wire stage2_c15_s_fa2;
    wire stage2_c15_c_fa2;
    wire stage2_c15_s_ha0;
    wire stage2_c15_c_ha0;
    wire stage2_c16_s_fa0;
    wire stage2_c16_c_fa0;
    wire stage2_c16_s_fa1;
    wire stage2_c16_c_fa1;
    wire stage2_c16_s_fa2;
    wire stage2_c16_c_fa2;
    wire stage2_c16_s_ha0;
    wire stage2_c16_c_ha0;
    wire stage2_c17_s_fa0;
    wire stage2_c17_c_fa0;
    wire stage2_c17_s_fa1;
    wire stage2_c17_c_fa1;
    wire stage2_c17_s_fa2;
    wire stage2_c17_c_fa2;
    wire stage2_c17_s_fa3;
    wire stage2_c17_c_fa3;
    wire stage2_c18_s_fa0;
    wire stage2_c18_c_fa0;
    wire stage2_c18_s_fa1;
    wire stage2_c18_c_fa1;
    wire stage2_c18_s_fa2;
    wire stage2_c18_c_fa2;
    wire stage2_c18_s_fa3;
    wire stage2_c18_c_fa3;
    wire stage2_c19_s_fa0;
    wire stage2_c19_c_fa0;
    wire stage2_c19_s_fa1;
    wire stage2_c19_c_fa1;
    wire stage2_c19_s_fa2;
    wire stage2_c19_c_fa2;
    wire stage2_c19_s_fa3;
    wire stage2_c19_c_fa3;
    wire stage2_c20_s_fa0;
    wire stage2_c20_c_fa0;
    wire stage2_c20_s_fa1;
    wire stage2_c20_c_fa1;
    wire stage2_c20_s_fa2;
    wire stage2_c20_c_fa2;
    wire stage2_c20_s_fa3;
    wire stage2_c20_c_fa3;
    wire stage2_c20_s_ha0;
    wire stage2_c20_c_ha0;
    wire stage2_c21_s_fa0;
    wire stage2_c21_c_fa0;
    wire stage2_c21_s_fa1;
    wire stage2_c21_c_fa1;
    wire stage2_c21_s_fa2;
    wire stage2_c21_c_fa2;
    wire stage2_c21_s_fa3;
    wire stage2_c21_c_fa3;
    wire stage2_c21_s_fa4;
    wire stage2_c21_c_fa4;
    wire stage2_c22_s_fa0;
    wire stage2_c22_c_fa0;
    wire stage2_c22_s_fa1;
    wire stage2_c22_c_fa1;
    wire stage2_c22_s_fa2;
    wire stage2_c22_c_fa2;
    wire stage2_c22_s_fa3;
    wire stage2_c22_c_fa3;
    wire stage2_c22_s_fa4;
    wire stage2_c22_c_fa4;
    wire stage2_c23_s_fa0;
    wire stage2_c23_c_fa0;
    wire stage2_c23_s_fa1;
    wire stage2_c23_c_fa1;
    wire stage2_c23_s_fa2;
    wire stage2_c23_c_fa2;
    wire stage2_c23_s_fa3;
    wire stage2_c23_c_fa3;
    wire stage2_c23_s_fa4;
    wire stage2_c23_c_fa4;
    wire stage2_c24_s_fa0;
    wire stage2_c24_c_fa0;
    wire stage2_c24_s_fa1;
    wire stage2_c24_c_fa1;
    wire stage2_c24_s_fa2;
    wire stage2_c24_c_fa2;
    wire stage2_c24_s_fa3;
    wire stage2_c24_c_fa3;
    wire stage2_c24_s_fa4;
    wire stage2_c24_c_fa4;
    wire stage2_c24_s_ha0;
    wire stage2_c24_c_ha0;
    wire stage2_c25_s_fa0;
    wire stage2_c25_c_fa0;
    wire stage2_c25_s_fa1;
    wire stage2_c25_c_fa1;
    wire stage2_c25_s_fa2;
    wire stage2_c25_c_fa2;
    wire stage2_c25_s_fa3;
    wire stage2_c25_c_fa3;
    wire stage2_c25_s_fa4;
    wire stage2_c25_c_fa4;
    wire stage2_c25_s_ha0;
    wire stage2_c25_c_ha0;
    wire stage2_c26_s_fa0;
    wire stage2_c26_c_fa0;
    wire stage2_c26_s_fa1;
    wire stage2_c26_c_fa1;
    wire stage2_c26_s_fa2;
    wire stage2_c26_c_fa2;
    wire stage2_c26_s_fa3;
    wire stage2_c26_c_fa3;
    wire stage2_c26_s_fa4;
    wire stage2_c26_c_fa4;
    wire stage2_c26_s_fa5;
    wire stage2_c26_c_fa5;
    wire stage2_c27_s_fa0;
    wire stage2_c27_c_fa0;
    wire stage2_c27_s_fa1;
    wire stage2_c27_c_fa1;
    wire stage2_c27_s_fa2;
    wire stage2_c27_c_fa2;
    wire stage2_c27_s_fa3;
    wire stage2_c27_c_fa3;
    wire stage2_c27_s_fa4;
    wire stage2_c27_c_fa4;
    wire stage2_c27_s_fa5;
    wire stage2_c27_c_fa5;
    wire stage2_c28_s_fa0;
    wire stage2_c28_c_fa0;
    wire stage2_c28_s_fa1;
    wire stage2_c28_c_fa1;
    wire stage2_c28_s_fa2;
    wire stage2_c28_c_fa2;
    wire stage2_c28_s_fa3;
    wire stage2_c28_c_fa3;
    wire stage2_c28_s_fa4;
    wire stage2_c28_c_fa4;
    wire stage2_c28_s_fa5;
    wire stage2_c28_c_fa5;
    wire stage2_c29_s_fa0;
    wire stage2_c29_c_fa0;
    wire stage2_c29_s_fa1;
    wire stage2_c29_c_fa1;
    wire stage2_c29_s_fa2;
    wire stage2_c29_c_fa2;
    wire stage2_c29_s_fa3;
    wire stage2_c29_c_fa3;
    wire stage2_c29_s_fa4;
    wire stage2_c29_c_fa4;
    wire stage2_c29_s_fa5;
    wire stage2_c29_c_fa5;
    wire stage2_c29_s_ha0;
    wire stage2_c29_c_ha0;
    wire stage2_c30_s_fa0;
    wire stage2_c30_c_fa0;
    wire stage2_c30_s_fa1;
    wire stage2_c30_c_fa1;
    wire stage2_c30_s_fa2;
    wire stage2_c30_c_fa2;
    wire stage2_c30_s_fa3;
    wire stage2_c30_c_fa3;
    wire stage2_c30_s_fa4;
    wire stage2_c30_c_fa4;
    wire stage2_c30_s_fa5;
    wire stage2_c30_c_fa5;
    wire stage2_c30_s_fa6;
    wire stage2_c30_c_fa6;
    wire stage2_c31_s_fa0;
    wire stage2_c31_c_fa0;
    wire stage2_c31_s_fa1;
    wire stage2_c31_c_fa1;
    wire stage2_c31_s_fa2;
    wire stage2_c31_c_fa2;
    wire stage2_c31_s_fa3;
    wire stage2_c31_c_fa3;
    wire stage2_c31_s_fa4;
    wire stage2_c31_c_fa4;
    wire stage2_c31_s_fa5;
    wire stage2_c31_c_fa5;
    wire stage2_c31_s_fa6;
    wire stage2_c31_c_fa6;
    wire stage2_c32_s_fa0;
    wire stage2_c32_c_fa0;
    wire stage2_c32_s_fa1;
    wire stage2_c32_c_fa1;
    wire stage2_c32_s_fa2;
    wire stage2_c32_c_fa2;
    wire stage2_c32_s_fa3;
    wire stage2_c32_c_fa3;
    wire stage2_c32_s_fa4;
    wire stage2_c32_c_fa4;
    wire stage2_c32_s_fa5;
    wire stage2_c32_c_fa5;
    wire stage2_c32_s_fa6;
    wire stage2_c32_c_fa6;
    wire stage2_c33_s_fa0;
    wire stage2_c33_c_fa0;
    wire stage2_c33_s_fa1;
    wire stage2_c33_c_fa1;
    wire stage2_c33_s_fa2;
    wire stage2_c33_c_fa2;
    wire stage2_c33_s_fa3;
    wire stage2_c33_c_fa3;
    wire stage2_c33_s_fa4;
    wire stage2_c33_c_fa4;
    wire stage2_c33_s_fa5;
    wire stage2_c33_c_fa5;
    wire stage2_c33_s_fa6;
    wire stage2_c33_c_fa6;
    wire stage2_c33_s_ha0;
    wire stage2_c33_c_ha0;
    wire stage2_c34_s_fa0;
    wire stage2_c34_c_fa0;
    wire stage2_c34_s_fa1;
    wire stage2_c34_c_fa1;
    wire stage2_c34_s_fa2;
    wire stage2_c34_c_fa2;
    wire stage2_c34_s_fa3;
    wire stage2_c34_c_fa3;
    wire stage2_c34_s_fa4;
    wire stage2_c34_c_fa4;
    wire stage2_c34_s_fa5;
    wire stage2_c34_c_fa5;
    wire stage2_c34_s_fa6;
    wire stage2_c34_c_fa6;
    wire stage2_c34_s_ha0;
    wire stage2_c34_c_ha0;
    wire stage2_c35_s_fa0;
    wire stage2_c35_c_fa0;
    wire stage2_c35_s_fa1;
    wire stage2_c35_c_fa1;
    wire stage2_c35_s_fa2;
    wire stage2_c35_c_fa2;
    wire stage2_c35_s_fa3;
    wire stage2_c35_c_fa3;
    wire stage2_c35_s_fa4;
    wire stage2_c35_c_fa4;
    wire stage2_c35_s_fa5;
    wire stage2_c35_c_fa5;
    wire stage2_c35_s_fa6;
    wire stage2_c35_c_fa6;
    wire stage2_c35_s_fa7;
    wire stage2_c35_c_fa7;
    wire stage2_c36_s_fa0;
    wire stage2_c36_c_fa0;
    wire stage2_c36_s_fa1;
    wire stage2_c36_c_fa1;
    wire stage2_c36_s_fa2;
    wire stage2_c36_c_fa2;
    wire stage2_c36_s_fa3;
    wire stage2_c36_c_fa3;
    wire stage2_c36_s_fa4;
    wire stage2_c36_c_fa4;
    wire stage2_c36_s_fa5;
    wire stage2_c36_c_fa5;
    wire stage2_c36_s_fa6;
    wire stage2_c36_c_fa6;
    wire stage2_c36_s_fa7;
    wire stage2_c36_c_fa7;
    wire stage2_c37_s_fa0;
    wire stage2_c37_c_fa0;
    wire stage2_c37_s_fa1;
    wire stage2_c37_c_fa1;
    wire stage2_c37_s_fa2;
    wire stage2_c37_c_fa2;
    wire stage2_c37_s_fa3;
    wire stage2_c37_c_fa3;
    wire stage2_c37_s_fa4;
    wire stage2_c37_c_fa4;
    wire stage2_c37_s_fa5;
    wire stage2_c37_c_fa5;
    wire stage2_c37_s_fa6;
    wire stage2_c37_c_fa6;
    wire stage2_c37_s_fa7;
    wire stage2_c37_c_fa7;
    wire stage2_c38_s_fa0;
    wire stage2_c38_c_fa0;
    wire stage2_c38_s_fa1;
    wire stage2_c38_c_fa1;
    wire stage2_c38_s_fa2;
    wire stage2_c38_c_fa2;
    wire stage2_c38_s_fa3;
    wire stage2_c38_c_fa3;
    wire stage2_c38_s_fa4;
    wire stage2_c38_c_fa4;
    wire stage2_c38_s_fa5;
    wire stage2_c38_c_fa5;
    wire stage2_c38_s_fa6;
    wire stage2_c38_c_fa6;
    wire stage2_c38_s_fa7;
    wire stage2_c38_c_fa7;
    wire stage2_c38_s_ha0;
    wire stage2_c38_c_ha0;
    wire stage2_c39_s_fa0;
    wire stage2_c39_c_fa0;
    wire stage2_c39_s_fa1;
    wire stage2_c39_c_fa1;
    wire stage2_c39_s_fa2;
    wire stage2_c39_c_fa2;
    wire stage2_c39_s_fa3;
    wire stage2_c39_c_fa3;
    wire stage2_c39_s_fa4;
    wire stage2_c39_c_fa4;
    wire stage2_c39_s_fa5;
    wire stage2_c39_c_fa5;
    wire stage2_c39_s_fa6;
    wire stage2_c39_c_fa6;
    wire stage2_c39_s_fa7;
    wire stage2_c39_c_fa7;
    wire stage2_c39_s_fa8;
    wire stage2_c39_c_fa8;
    wire stage2_c40_s_fa0;
    wire stage2_c40_c_fa0;
    wire stage2_c40_s_fa1;
    wire stage2_c40_c_fa1;
    wire stage2_c40_s_fa2;
    wire stage2_c40_c_fa2;
    wire stage2_c40_s_fa3;
    wire stage2_c40_c_fa3;
    wire stage2_c40_s_fa4;
    wire stage2_c40_c_fa4;
    wire stage2_c40_s_fa5;
    wire stage2_c40_c_fa5;
    wire stage2_c40_s_fa6;
    wire stage2_c40_c_fa6;
    wire stage2_c40_s_fa7;
    wire stage2_c40_c_fa7;
    wire stage2_c40_s_fa8;
    wire stage2_c40_c_fa8;
    wire stage2_c41_s_fa0;
    wire stage2_c41_c_fa0;
    wire stage2_c41_s_fa1;
    wire stage2_c41_c_fa1;
    wire stage2_c41_s_fa2;
    wire stage2_c41_c_fa2;
    wire stage2_c41_s_fa3;
    wire stage2_c41_c_fa3;
    wire stage2_c41_s_fa4;
    wire stage2_c41_c_fa4;
    wire stage2_c41_s_fa5;
    wire stage2_c41_c_fa5;
    wire stage2_c41_s_fa6;
    wire stage2_c41_c_fa6;
    wire stage2_c41_s_fa7;
    wire stage2_c41_c_fa7;
    wire stage2_c41_s_fa8;
    wire stage2_c41_c_fa8;
    wire stage2_c42_s_fa0;
    wire stage2_c42_c_fa0;
    wire stage2_c42_s_fa1;
    wire stage2_c42_c_fa1;
    wire stage2_c42_s_fa2;
    wire stage2_c42_c_fa2;
    wire stage2_c42_s_fa3;
    wire stage2_c42_c_fa3;
    wire stage2_c42_s_fa4;
    wire stage2_c42_c_fa4;
    wire stage2_c42_s_fa5;
    wire stage2_c42_c_fa5;
    wire stage2_c42_s_fa6;
    wire stage2_c42_c_fa6;
    wire stage2_c42_s_fa7;
    wire stage2_c42_c_fa7;
    wire stage2_c42_s_fa8;
    wire stage2_c42_c_fa8;
    wire stage2_c43_s_fa0;
    wire stage2_c43_c_fa0;
    wire stage2_c43_s_fa1;
    wire stage2_c43_c_fa1;
    wire stage2_c43_s_fa2;
    wire stage2_c43_c_fa2;
    wire stage2_c43_s_fa3;
    wire stage2_c43_c_fa3;
    wire stage2_c43_s_fa4;
    wire stage2_c43_c_fa4;
    wire stage2_c43_s_fa5;
    wire stage2_c43_c_fa5;
    wire stage2_c43_s_fa6;
    wire stage2_c43_c_fa6;
    wire stage2_c43_s_fa7;
    wire stage2_c43_c_fa7;
    wire stage2_c43_s_fa8;
    wire stage2_c43_c_fa8;
    wire stage2_c44_s_fa0;
    wire stage2_c44_c_fa0;
    wire stage2_c44_s_fa1;
    wire stage2_c44_c_fa1;
    wire stage2_c44_s_fa2;
    wire stage2_c44_c_fa2;
    wire stage2_c44_s_fa3;
    wire stage2_c44_c_fa3;
    wire stage2_c44_s_fa4;
    wire stage2_c44_c_fa4;
    wire stage2_c44_s_fa5;
    wire stage2_c44_c_fa5;
    wire stage2_c44_s_fa6;
    wire stage2_c44_c_fa6;
    wire stage2_c44_s_fa7;
    wire stage2_c44_c_fa7;
    wire stage2_c44_s_fa8;
    wire stage2_c44_c_fa8;
    wire stage2_c45_s_fa0;
    wire stage2_c45_c_fa0;
    wire stage2_c45_s_fa1;
    wire stage2_c45_c_fa1;
    wire stage2_c45_s_fa2;
    wire stage2_c45_c_fa2;
    wire stage2_c45_s_fa3;
    wire stage2_c45_c_fa3;
    wire stage2_c45_s_fa4;
    wire stage2_c45_c_fa4;
    wire stage2_c45_s_fa5;
    wire stage2_c45_c_fa5;
    wire stage2_c45_s_fa6;
    wire stage2_c45_c_fa6;
    wire stage2_c45_s_fa7;
    wire stage2_c45_c_fa7;
    wire stage2_c45_s_fa8;
    wire stage2_c45_c_fa8;
    wire stage2_c46_s_fa0;
    wire stage2_c46_c_fa0;
    wire stage2_c46_s_fa1;
    wire stage2_c46_c_fa1;
    wire stage2_c46_s_fa2;
    wire stage2_c46_c_fa2;
    wire stage2_c46_s_fa3;
    wire stage2_c46_c_fa3;
    wire stage2_c46_s_fa4;
    wire stage2_c46_c_fa4;
    wire stage2_c46_s_fa5;
    wire stage2_c46_c_fa5;
    wire stage2_c46_s_fa6;
    wire stage2_c46_c_fa6;
    wire stage2_c46_s_fa7;
    wire stage2_c46_c_fa7;
    wire stage2_c46_s_fa8;
    wire stage2_c46_c_fa8;
    wire stage2_c47_s_fa0;
    wire stage2_c47_c_fa0;
    wire stage2_c47_s_fa1;
    wire stage2_c47_c_fa1;
    wire stage2_c47_s_fa2;
    wire stage2_c47_c_fa2;
    wire stage2_c47_s_fa3;
    wire stage2_c47_c_fa3;
    wire stage2_c47_s_fa4;
    wire stage2_c47_c_fa4;
    wire stage2_c47_s_fa5;
    wire stage2_c47_c_fa5;
    wire stage2_c47_s_fa6;
    wire stage2_c47_c_fa6;
    wire stage2_c47_s_fa7;
    wire stage2_c47_c_fa7;
    wire stage2_c47_s_fa8;
    wire stage2_c47_c_fa8;
    wire stage2_c48_s_fa0;
    wire stage2_c48_c_fa0;
    wire stage2_c48_s_fa1;
    wire stage2_c48_c_fa1;
    wire stage2_c48_s_fa2;
    wire stage2_c48_c_fa2;
    wire stage2_c48_s_fa3;
    wire stage2_c48_c_fa3;
    wire stage2_c48_s_fa4;
    wire stage2_c48_c_fa4;
    wire stage2_c48_s_fa5;
    wire stage2_c48_c_fa5;
    wire stage2_c48_s_fa6;
    wire stage2_c48_c_fa6;
    wire stage2_c48_s_fa7;
    wire stage2_c48_c_fa7;
    wire stage2_c48_s_fa8;
    wire stage2_c48_c_fa8;
    wire stage2_c49_s_fa0;
    wire stage2_c49_c_fa0;
    wire stage2_c49_s_fa1;
    wire stage2_c49_c_fa1;
    wire stage2_c49_s_fa2;
    wire stage2_c49_c_fa2;
    wire stage2_c49_s_fa3;
    wire stage2_c49_c_fa3;
    wire stage2_c49_s_fa4;
    wire stage2_c49_c_fa4;
    wire stage2_c49_s_fa5;
    wire stage2_c49_c_fa5;
    wire stage2_c49_s_fa6;
    wire stage2_c49_c_fa6;
    wire stage2_c49_s_fa7;
    wire stage2_c49_c_fa7;
    wire stage2_c49_s_fa8;
    wire stage2_c49_c_fa8;
    wire stage2_c50_s_fa0;
    wire stage2_c50_c_fa0;
    wire stage2_c50_s_fa1;
    wire stage2_c50_c_fa1;
    wire stage2_c50_s_fa2;
    wire stage2_c50_c_fa2;
    wire stage2_c50_s_fa3;
    wire stage2_c50_c_fa3;
    wire stage2_c50_s_fa4;
    wire stage2_c50_c_fa4;
    wire stage2_c50_s_fa5;
    wire stage2_c50_c_fa5;
    wire stage2_c50_s_fa6;
    wire stage2_c50_c_fa6;
    wire stage2_c50_s_fa7;
    wire stage2_c50_c_fa7;
    wire stage2_c50_s_fa8;
    wire stage2_c50_c_fa8;
    wire stage2_c51_s_fa0;
    wire stage2_c51_c_fa0;
    wire stage2_c51_s_fa1;
    wire stage2_c51_c_fa1;
    wire stage2_c51_s_fa2;
    wire stage2_c51_c_fa2;
    wire stage2_c51_s_fa3;
    wire stage2_c51_c_fa3;
    wire stage2_c51_s_fa4;
    wire stage2_c51_c_fa4;
    wire stage2_c51_s_fa5;
    wire stage2_c51_c_fa5;
    wire stage2_c51_s_fa6;
    wire stage2_c51_c_fa6;
    wire stage2_c51_s_fa7;
    wire stage2_c51_c_fa7;
    wire stage2_c51_s_fa8;
    wire stage2_c51_c_fa8;
    wire stage2_c52_s_fa0;
    wire stage2_c52_c_fa0;
    wire stage2_c52_s_fa1;
    wire stage2_c52_c_fa1;
    wire stage2_c52_s_fa2;
    wire stage2_c52_c_fa2;
    wire stage2_c52_s_fa3;
    wire stage2_c52_c_fa3;
    wire stage2_c52_s_fa4;
    wire stage2_c52_c_fa4;
    wire stage2_c52_s_fa5;
    wire stage2_c52_c_fa5;
    wire stage2_c52_s_fa6;
    wire stage2_c52_c_fa6;
    wire stage2_c52_s_fa7;
    wire stage2_c52_c_fa7;
    wire stage2_c52_s_fa8;
    wire stage2_c52_c_fa8;
    wire stage2_c53_s_fa0;
    wire stage2_c53_c_fa0;
    wire stage2_c53_s_fa1;
    wire stage2_c53_c_fa1;
    wire stage2_c53_s_fa2;
    wire stage2_c53_c_fa2;
    wire stage2_c53_s_fa3;
    wire stage2_c53_c_fa3;
    wire stage2_c53_s_fa4;
    wire stage2_c53_c_fa4;
    wire stage2_c53_s_fa5;
    wire stage2_c53_c_fa5;
    wire stage2_c53_s_fa6;
    wire stage2_c53_c_fa6;
    wire stage2_c53_s_fa7;
    wire stage2_c53_c_fa7;
    wire stage2_c53_s_fa8;
    wire stage2_c53_c_fa8;
    wire stage2_c54_s_fa0;
    wire stage2_c54_c_fa0;
    wire stage2_c54_s_fa1;
    wire stage2_c54_c_fa1;
    wire stage2_c54_s_fa2;
    wire stage2_c54_c_fa2;
    wire stage2_c54_s_fa3;
    wire stage2_c54_c_fa3;
    wire stage2_c54_s_fa4;
    wire stage2_c54_c_fa4;
    wire stage2_c54_s_fa5;
    wire stage2_c54_c_fa5;
    wire stage2_c54_s_fa6;
    wire stage2_c54_c_fa6;
    wire stage2_c54_s_fa7;
    wire stage2_c54_c_fa7;
    wire stage2_c54_s_fa8;
    wire stage2_c54_c_fa8;
    wire stage2_c55_s_fa0;
    wire stage2_c55_c_fa0;
    wire stage2_c55_s_fa1;
    wire stage2_c55_c_fa1;
    wire stage2_c55_s_fa2;
    wire stage2_c55_c_fa2;
    wire stage2_c55_s_fa3;
    wire stage2_c55_c_fa3;
    wire stage2_c55_s_fa4;
    wire stage2_c55_c_fa4;
    wire stage2_c55_s_fa5;
    wire stage2_c55_c_fa5;
    wire stage2_c55_s_fa6;
    wire stage2_c55_c_fa6;
    wire stage2_c55_s_fa7;
    wire stage2_c55_c_fa7;
    wire stage2_c55_s_fa8;
    wire stage2_c55_c_fa8;
    wire stage2_c56_s_fa0;
    wire stage2_c56_c_fa0;
    wire stage2_c56_s_fa1;
    wire stage2_c56_c_fa1;
    wire stage2_c56_s_fa2;
    wire stage2_c56_c_fa2;
    wire stage2_c56_s_fa3;
    wire stage2_c56_c_fa3;
    wire stage2_c56_s_fa4;
    wire stage2_c56_c_fa4;
    wire stage2_c56_s_fa5;
    wire stage2_c56_c_fa5;
    wire stage2_c56_s_fa6;
    wire stage2_c56_c_fa6;
    wire stage2_c56_s_fa7;
    wire stage2_c56_c_fa7;
    wire stage2_c56_s_fa8;
    wire stage2_c56_c_fa8;
    wire stage2_c57_s_fa0;
    wire stage2_c57_c_fa0;
    wire stage2_c57_s_fa1;
    wire stage2_c57_c_fa1;
    wire stage2_c57_s_fa2;
    wire stage2_c57_c_fa2;
    wire stage2_c57_s_fa3;
    wire stage2_c57_c_fa3;
    wire stage2_c57_s_fa4;
    wire stage2_c57_c_fa4;
    wire stage2_c57_s_fa5;
    wire stage2_c57_c_fa5;
    wire stage2_c57_s_fa6;
    wire stage2_c57_c_fa6;
    wire stage2_c57_s_fa7;
    wire stage2_c57_c_fa7;
    wire stage2_c57_s_fa8;
    wire stage2_c57_c_fa8;
    wire stage2_c58_s_fa0;
    wire stage2_c58_c_fa0;
    wire stage2_c58_s_fa1;
    wire stage2_c58_c_fa1;
    wire stage2_c58_s_fa2;
    wire stage2_c58_c_fa2;
    wire stage2_c58_s_fa3;
    wire stage2_c58_c_fa3;
    wire stage2_c58_s_fa4;
    wire stage2_c58_c_fa4;
    wire stage2_c58_s_fa5;
    wire stage2_c58_c_fa5;
    wire stage2_c58_s_fa6;
    wire stage2_c58_c_fa6;
    wire stage2_c58_s_fa7;
    wire stage2_c58_c_fa7;
    wire stage2_c58_s_fa8;
    wire stage2_c58_c_fa8;
    wire stage2_c59_s_fa0;
    wire stage2_c59_c_fa0;
    wire stage2_c59_s_fa1;
    wire stage2_c59_c_fa1;
    wire stage2_c59_s_fa2;
    wire stage2_c59_c_fa2;
    wire stage2_c59_s_fa3;
    wire stage2_c59_c_fa3;
    wire stage2_c59_s_fa4;
    wire stage2_c59_c_fa4;
    wire stage2_c59_s_fa5;
    wire stage2_c59_c_fa5;
    wire stage2_c59_s_fa6;
    wire stage2_c59_c_fa6;
    wire stage2_c59_s_fa7;
    wire stage2_c59_c_fa7;
    wire stage2_c59_s_fa8;
    wire stage2_c59_c_fa8;
    wire stage2_c60_s_fa0;
    wire stage2_c60_c_fa0;
    wire stage2_c60_s_fa1;
    wire stage2_c60_c_fa1;
    wire stage2_c60_s_fa2;
    wire stage2_c60_c_fa2;
    wire stage2_c60_s_fa3;
    wire stage2_c60_c_fa3;
    wire stage2_c60_s_fa4;
    wire stage2_c60_c_fa4;
    wire stage2_c60_s_fa5;
    wire stage2_c60_c_fa5;
    wire stage2_c60_s_fa6;
    wire stage2_c60_c_fa6;
    wire stage2_c60_s_fa7;
    wire stage2_c60_c_fa7;
    wire stage2_c60_s_fa8;
    wire stage2_c60_c_fa8;
    wire stage2_c61_s_fa0;
    wire stage2_c61_c_fa0;
    wire stage2_c61_s_fa1;
    wire stage2_c61_c_fa1;
    wire stage2_c61_s_fa2;
    wire stage2_c61_c_fa2;
    wire stage2_c61_s_fa3;
    wire stage2_c61_c_fa3;
    wire stage2_c61_s_fa4;
    wire stage2_c61_c_fa4;
    wire stage2_c61_s_fa5;
    wire stage2_c61_c_fa5;
    wire stage2_c61_s_fa6;
    wire stage2_c61_c_fa6;
    wire stage2_c61_s_fa7;
    wire stage2_c61_c_fa7;
    wire stage2_c61_s_fa8;
    wire stage2_c61_c_fa8;
    wire stage2_c62_s_fa0;
    wire stage2_c62_c_fa0;
    wire stage2_c62_s_fa1;
    wire stage2_c62_c_fa1;
    wire stage2_c62_s_fa2;
    wire stage2_c62_c_fa2;
    wire stage2_c62_s_fa3;
    wire stage2_c62_c_fa3;
    wire stage2_c62_s_fa4;
    wire stage2_c62_c_fa4;
    wire stage2_c62_s_fa5;
    wire stage2_c62_c_fa5;
    wire stage2_c62_s_fa6;
    wire stage2_c62_c_fa6;
    wire stage2_c62_s_fa7;
    wire stage2_c62_c_fa7;
    wire stage2_c62_s_fa8;
    wire stage2_c62_c_fa8;
    wire stage2_c63_s_fa0;
    wire stage2_c63_c_fa0;
    wire stage2_c63_s_fa1;
    wire stage2_c63_c_fa1;
    wire stage2_c63_s_fa2;
    wire stage2_c63_c_fa2;
    wire stage2_c63_s_fa3;
    wire stage2_c63_c_fa3;
    wire stage2_c63_s_fa4;
    wire stage2_c63_c_fa4;
    wire stage2_c63_s_fa5;
    wire stage2_c63_c_fa5;
    wire stage2_c63_s_fa6;
    wire stage2_c63_c_fa6;
    wire stage2_c63_s_fa7;
    wire stage2_c63_c_fa7;
    wire stage2_c63_s_fa8;
    wire stage2_c63_c_fa8;
    wire stage2_c64_s_fa0;
    wire stage2_c64_c_fa0;
    wire stage2_c64_s_fa1;
    wire stage2_c64_c_fa1;
    wire stage2_c64_s_fa2;
    wire stage2_c64_c_fa2;
    wire stage2_c64_s_fa3;
    wire stage2_c64_c_fa3;
    wire stage2_c64_s_fa4;
    wire stage2_c64_c_fa4;
    wire stage2_c64_s_fa5;
    wire stage2_c64_c_fa5;
    wire stage2_c64_s_fa6;
    wire stage2_c64_c_fa6;
    wire stage2_c64_s_fa7;
    wire stage2_c64_c_fa7;
    wire stage2_c64_s_fa8;
    wire stage2_c64_c_fa8;
    wire stage2_c65_s_fa0;
    wire stage2_c65_c_fa0;
    wire stage2_c65_s_fa1;
    wire stage2_c65_c_fa1;
    wire stage2_c65_s_fa2;
    wire stage2_c65_c_fa2;
    wire stage2_c65_s_fa3;
    wire stage2_c65_c_fa3;
    wire stage2_c65_s_fa4;
    wire stage2_c65_c_fa4;
    wire stage2_c65_s_fa5;
    wire stage2_c65_c_fa5;
    wire stage2_c65_s_fa6;
    wire stage2_c65_c_fa6;
    wire stage2_c65_s_fa7;
    wire stage2_c65_c_fa7;
    wire stage2_c65_s_fa8;
    wire stage2_c65_c_fa8;
    wire stage2_c66_s_fa0;
    wire stage2_c66_c_fa0;
    wire stage2_c66_s_fa1;
    wire stage2_c66_c_fa1;
    wire stage2_c66_s_fa2;
    wire stage2_c66_c_fa2;
    wire stage2_c66_s_fa3;
    wire stage2_c66_c_fa3;
    wire stage2_c66_s_fa4;
    wire stage2_c66_c_fa4;
    wire stage2_c66_s_fa5;
    wire stage2_c66_c_fa5;
    wire stage2_c66_s_fa6;
    wire stage2_c66_c_fa6;
    wire stage2_c66_s_fa7;
    wire stage2_c66_c_fa7;
    wire stage2_c66_s_fa8;
    wire stage2_c66_c_fa8;
    wire stage2_c67_s_fa0;
    wire stage2_c67_c_fa0;
    wire stage2_c67_s_fa1;
    wire stage2_c67_c_fa1;
    wire stage2_c67_s_fa2;
    wire stage2_c67_c_fa2;
    wire stage2_c67_s_fa3;
    wire stage2_c67_c_fa3;
    wire stage2_c67_s_fa4;
    wire stage2_c67_c_fa4;
    wire stage2_c67_s_fa5;
    wire stage2_c67_c_fa5;
    wire stage2_c67_s_fa6;
    wire stage2_c67_c_fa6;
    wire stage2_c67_s_fa7;
    wire stage2_c67_c_fa7;
    wire stage2_c67_s_fa8;
    wire stage2_c67_c_fa8;
    wire stage2_c68_s_fa0;
    wire stage2_c68_c_fa0;
    wire stage2_c68_s_fa1;
    wire stage2_c68_c_fa1;
    wire stage2_c68_s_fa2;
    wire stage2_c68_c_fa2;
    wire stage2_c68_s_fa3;
    wire stage2_c68_c_fa3;
    wire stage2_c68_s_fa4;
    wire stage2_c68_c_fa4;
    wire stage2_c68_s_fa5;
    wire stage2_c68_c_fa5;
    wire stage2_c68_s_fa6;
    wire stage2_c68_c_fa6;
    wire stage2_c68_s_fa7;
    wire stage2_c68_c_fa7;
    wire stage2_c68_s_fa8;
    wire stage2_c68_c_fa8;
    wire stage2_c69_s_fa0;
    wire stage2_c69_c_fa0;
    wire stage2_c69_s_fa1;
    wire stage2_c69_c_fa1;
    wire stage2_c69_s_fa2;
    wire stage2_c69_c_fa2;
    wire stage2_c69_s_fa3;
    wire stage2_c69_c_fa3;
    wire stage2_c69_s_fa4;
    wire stage2_c69_c_fa4;
    wire stage2_c69_s_fa5;
    wire stage2_c69_c_fa5;
    wire stage2_c69_s_fa6;
    wire stage2_c69_c_fa6;
    wire stage2_c69_s_fa7;
    wire stage2_c69_c_fa7;
    wire stage2_c69_s_fa8;
    wire stage2_c69_c_fa8;
    wire stage2_c70_s_fa0;
    wire stage2_c70_c_fa0;
    wire stage2_c70_s_fa1;
    wire stage2_c70_c_fa1;
    wire stage2_c70_s_fa2;
    wire stage2_c70_c_fa2;
    wire stage2_c70_s_fa3;
    wire stage2_c70_c_fa3;
    wire stage2_c70_s_fa4;
    wire stage2_c70_c_fa4;
    wire stage2_c70_s_fa5;
    wire stage2_c70_c_fa5;
    wire stage2_c70_s_fa6;
    wire stage2_c70_c_fa6;
    wire stage2_c70_s_fa7;
    wire stage2_c70_c_fa7;
    wire stage2_c70_s_fa8;
    wire stage2_c70_c_fa8;
    wire stage2_c71_s_fa0;
    wire stage2_c71_c_fa0;
    wire stage2_c71_s_fa1;
    wire stage2_c71_c_fa1;
    wire stage2_c71_s_fa2;
    wire stage2_c71_c_fa2;
    wire stage2_c71_s_fa3;
    wire stage2_c71_c_fa3;
    wire stage2_c71_s_fa4;
    wire stage2_c71_c_fa4;
    wire stage2_c71_s_fa5;
    wire stage2_c71_c_fa5;
    wire stage2_c71_s_fa6;
    wire stage2_c71_c_fa6;
    wire stage2_c71_s_fa7;
    wire stage2_c71_c_fa7;
    wire stage2_c71_s_fa8;
    wire stage2_c71_c_fa8;
    wire stage2_c72_s_fa0;
    wire stage2_c72_c_fa0;
    wire stage2_c72_s_fa1;
    wire stage2_c72_c_fa1;
    wire stage2_c72_s_fa2;
    wire stage2_c72_c_fa2;
    wire stage2_c72_s_fa3;
    wire stage2_c72_c_fa3;
    wire stage2_c72_s_fa4;
    wire stage2_c72_c_fa4;
    wire stage2_c72_s_fa5;
    wire stage2_c72_c_fa5;
    wire stage2_c72_s_fa6;
    wire stage2_c72_c_fa6;
    wire stage2_c72_s_fa7;
    wire stage2_c72_c_fa7;
    wire stage2_c72_s_fa8;
    wire stage2_c72_c_fa8;
    wire stage2_c73_s_fa0;
    wire stage2_c73_c_fa0;
    wire stage2_c73_s_fa1;
    wire stage2_c73_c_fa1;
    wire stage2_c73_s_fa2;
    wire stage2_c73_c_fa2;
    wire stage2_c73_s_fa3;
    wire stage2_c73_c_fa3;
    wire stage2_c73_s_fa4;
    wire stage2_c73_c_fa4;
    wire stage2_c73_s_fa5;
    wire stage2_c73_c_fa5;
    wire stage2_c73_s_fa6;
    wire stage2_c73_c_fa6;
    wire stage2_c73_s_fa7;
    wire stage2_c73_c_fa7;
    wire stage2_c73_s_ha0;
    wire stage2_c73_c_ha0;
    wire stage2_c74_s_fa0;
    wire stage2_c74_c_fa0;
    wire stage2_c74_s_fa1;
    wire stage2_c74_c_fa1;
    wire stage2_c74_s_fa2;
    wire stage2_c74_c_fa2;
    wire stage2_c74_s_fa3;
    wire stage2_c74_c_fa3;
    wire stage2_c74_s_fa4;
    wire stage2_c74_c_fa4;
    wire stage2_c74_s_fa5;
    wire stage2_c74_c_fa5;
    wire stage2_c74_s_fa6;
    wire stage2_c74_c_fa6;
    wire stage2_c74_s_fa7;
    wire stage2_c74_c_fa7;
    wire stage2_c74_s_ha0;
    wire stage2_c74_c_ha0;
    wire stage2_c75_s_fa0;
    wire stage2_c75_c_fa0;
    wire stage2_c75_s_fa1;
    wire stage2_c75_c_fa1;
    wire stage2_c75_s_fa2;
    wire stage2_c75_c_fa2;
    wire stage2_c75_s_fa3;
    wire stage2_c75_c_fa3;
    wire stage2_c75_s_fa4;
    wire stage2_c75_c_fa4;
    wire stage2_c75_s_fa5;
    wire stage2_c75_c_fa5;
    wire stage2_c75_s_fa6;
    wire stage2_c75_c_fa6;
    wire stage2_c75_s_fa7;
    wire stage2_c75_c_fa7;
    wire stage2_c75_s_ha0;
    wire stage2_c75_c_ha0;
    wire stage2_c76_s_fa0;
    wire stage2_c76_c_fa0;
    wire stage2_c76_s_fa1;
    wire stage2_c76_c_fa1;
    wire stage2_c76_s_fa2;
    wire stage2_c76_c_fa2;
    wire stage2_c76_s_fa3;
    wire stage2_c76_c_fa3;
    wire stage2_c76_s_fa4;
    wire stage2_c76_c_fa4;
    wire stage2_c76_s_fa5;
    wire stage2_c76_c_fa5;
    wire stage2_c76_s_fa6;
    wire stage2_c76_c_fa6;
    wire stage2_c76_s_fa7;
    wire stage2_c76_c_fa7;
    wire stage2_c77_s_fa0;
    wire stage2_c77_c_fa0;
    wire stage2_c77_s_fa1;
    wire stage2_c77_c_fa1;
    wire stage2_c77_s_fa2;
    wire stage2_c77_c_fa2;
    wire stage2_c77_s_fa3;
    wire stage2_c77_c_fa3;
    wire stage2_c77_s_fa4;
    wire stage2_c77_c_fa4;
    wire stage2_c77_s_fa5;
    wire stage2_c77_c_fa5;
    wire stage2_c77_s_fa6;
    wire stage2_c77_c_fa6;
    wire stage2_c77_s_fa7;
    wire stage2_c77_c_fa7;
    wire stage2_c78_s_fa0;
    wire stage2_c78_c_fa0;
    wire stage2_c78_s_fa1;
    wire stage2_c78_c_fa1;
    wire stage2_c78_s_fa2;
    wire stage2_c78_c_fa2;
    wire stage2_c78_s_fa3;
    wire stage2_c78_c_fa3;
    wire stage2_c78_s_fa4;
    wire stage2_c78_c_fa4;
    wire stage2_c78_s_fa5;
    wire stage2_c78_c_fa5;
    wire stage2_c78_s_fa6;
    wire stage2_c78_c_fa6;
    wire stage2_c78_s_fa7;
    wire stage2_c78_c_fa7;
    wire stage2_c79_s_fa0;
    wire stage2_c79_c_fa0;
    wire stage2_c79_s_fa1;
    wire stage2_c79_c_fa1;
    wire stage2_c79_s_fa2;
    wire stage2_c79_c_fa2;
    wire stage2_c79_s_fa3;
    wire stage2_c79_c_fa3;
    wire stage2_c79_s_fa4;
    wire stage2_c79_c_fa4;
    wire stage2_c79_s_fa5;
    wire stage2_c79_c_fa5;
    wire stage2_c79_s_fa6;
    wire stage2_c79_c_fa6;
    wire stage2_c80_s_fa0;
    wire stage2_c80_c_fa0;
    wire stage2_c80_s_fa1;
    wire stage2_c80_c_fa1;
    wire stage2_c80_s_fa2;
    wire stage2_c80_c_fa2;
    wire stage2_c80_s_fa3;
    wire stage2_c80_c_fa3;
    wire stage2_c80_s_fa4;
    wire stage2_c80_c_fa4;
    wire stage2_c80_s_fa5;
    wire stage2_c80_c_fa5;
    wire stage2_c80_s_fa6;
    wire stage2_c80_c_fa6;
    wire stage2_c81_s_fa0;
    wire stage2_c81_c_fa0;
    wire stage2_c81_s_fa1;
    wire stage2_c81_c_fa1;
    wire stage2_c81_s_fa2;
    wire stage2_c81_c_fa2;
    wire stage2_c81_s_fa3;
    wire stage2_c81_c_fa3;
    wire stage2_c81_s_fa4;
    wire stage2_c81_c_fa4;
    wire stage2_c81_s_fa5;
    wire stage2_c81_c_fa5;
    wire stage2_c81_s_fa6;
    wire stage2_c81_c_fa6;
    wire stage2_c82_s_fa0;
    wire stage2_c82_c_fa0;
    wire stage2_c82_s_fa1;
    wire stage2_c82_c_fa1;
    wire stage2_c82_s_fa2;
    wire stage2_c82_c_fa2;
    wire stage2_c82_s_fa3;
    wire stage2_c82_c_fa3;
    wire stage2_c82_s_fa4;
    wire stage2_c82_c_fa4;
    wire stage2_c82_s_fa5;
    wire stage2_c82_c_fa5;
    wire stage2_c82_s_ha0;
    wire stage2_c82_c_ha0;
    wire stage2_c83_s_fa0;
    wire stage2_c83_c_fa0;
    wire stage2_c83_s_fa1;
    wire stage2_c83_c_fa1;
    wire stage2_c83_s_fa2;
    wire stage2_c83_c_fa2;
    wire stage2_c83_s_fa3;
    wire stage2_c83_c_fa3;
    wire stage2_c83_s_fa4;
    wire stage2_c83_c_fa4;
    wire stage2_c83_s_fa5;
    wire stage2_c83_c_fa5;
    wire stage2_c83_s_ha0;
    wire stage2_c83_c_ha0;
    wire stage2_c84_s_fa0;
    wire stage2_c84_c_fa0;
    wire stage2_c84_s_fa1;
    wire stage2_c84_c_fa1;
    wire stage2_c84_s_fa2;
    wire stage2_c84_c_fa2;
    wire stage2_c84_s_fa3;
    wire stage2_c84_c_fa3;
    wire stage2_c84_s_fa4;
    wire stage2_c84_c_fa4;
    wire stage2_c84_s_fa5;
    wire stage2_c84_c_fa5;
    wire stage2_c84_s_ha0;
    wire stage2_c84_c_ha0;
    wire stage2_c85_s_fa0;
    wire stage2_c85_c_fa0;
    wire stage2_c85_s_fa1;
    wire stage2_c85_c_fa1;
    wire stage2_c85_s_fa2;
    wire stage2_c85_c_fa2;
    wire stage2_c85_s_fa3;
    wire stage2_c85_c_fa3;
    wire stage2_c85_s_fa4;
    wire stage2_c85_c_fa4;
    wire stage2_c85_s_fa5;
    wire stage2_c85_c_fa5;
    wire stage2_c86_s_fa0;
    wire stage2_c86_c_fa0;
    wire stage2_c86_s_fa1;
    wire stage2_c86_c_fa1;
    wire stage2_c86_s_fa2;
    wire stage2_c86_c_fa2;
    wire stage2_c86_s_fa3;
    wire stage2_c86_c_fa3;
    wire stage2_c86_s_fa4;
    wire stage2_c86_c_fa4;
    wire stage2_c86_s_fa5;
    wire stage2_c86_c_fa5;
    wire stage2_c87_s_fa0;
    wire stage2_c87_c_fa0;
    wire stage2_c87_s_fa1;
    wire stage2_c87_c_fa1;
    wire stage2_c87_s_fa2;
    wire stage2_c87_c_fa2;
    wire stage2_c87_s_fa3;
    wire stage2_c87_c_fa3;
    wire stage2_c87_s_fa4;
    wire stage2_c87_c_fa4;
    wire stage2_c87_s_fa5;
    wire stage2_c87_c_fa5;
    wire stage2_c88_s_fa0;
    wire stage2_c88_c_fa0;
    wire stage2_c88_s_fa1;
    wire stage2_c88_c_fa1;
    wire stage2_c88_s_fa2;
    wire stage2_c88_c_fa2;
    wire stage2_c88_s_fa3;
    wire stage2_c88_c_fa3;
    wire stage2_c88_s_fa4;
    wire stage2_c88_c_fa4;
    wire stage2_c89_s_fa0;
    wire stage2_c89_c_fa0;
    wire stage2_c89_s_fa1;
    wire stage2_c89_c_fa1;
    wire stage2_c89_s_fa2;
    wire stage2_c89_c_fa2;
    wire stage2_c89_s_fa3;
    wire stage2_c89_c_fa3;
    wire stage2_c89_s_fa4;
    wire stage2_c89_c_fa4;
    wire stage2_c90_s_fa0;
    wire stage2_c90_c_fa0;
    wire stage2_c90_s_fa1;
    wire stage2_c90_c_fa1;
    wire stage2_c90_s_fa2;
    wire stage2_c90_c_fa2;
    wire stage2_c90_s_fa3;
    wire stage2_c90_c_fa3;
    wire stage2_c90_s_fa4;
    wire stage2_c90_c_fa4;
    wire stage2_c91_s_fa0;
    wire stage2_c91_c_fa0;
    wire stage2_c91_s_fa1;
    wire stage2_c91_c_fa1;
    wire stage2_c91_s_fa2;
    wire stage2_c91_c_fa2;
    wire stage2_c91_s_fa3;
    wire stage2_c91_c_fa3;
    wire stage2_c91_s_ha0;
    wire stage2_c91_c_ha0;
    wire stage2_c92_s_fa0;
    wire stage2_c92_c_fa0;
    wire stage2_c92_s_fa1;
    wire stage2_c92_c_fa1;
    wire stage2_c92_s_fa2;
    wire stage2_c92_c_fa2;
    wire stage2_c92_s_fa3;
    wire stage2_c92_c_fa3;
    wire stage2_c92_s_ha0;
    wire stage2_c92_c_ha0;
    wire stage2_c93_s_fa0;
    wire stage2_c93_c_fa0;
    wire stage2_c93_s_fa1;
    wire stage2_c93_c_fa1;
    wire stage2_c93_s_fa2;
    wire stage2_c93_c_fa2;
    wire stage2_c93_s_fa3;
    wire stage2_c93_c_fa3;
    wire stage2_c93_s_ha0;
    wire stage2_c93_c_ha0;
    wire stage2_c94_s_fa0;
    wire stage2_c94_c_fa0;
    wire stage2_c94_s_fa1;
    wire stage2_c94_c_fa1;
    wire stage2_c94_s_fa2;
    wire stage2_c94_c_fa2;
    wire stage2_c94_s_fa3;
    wire stage2_c94_c_fa3;
    wire stage2_c95_s_fa0;
    wire stage2_c95_c_fa0;
    wire stage2_c95_s_fa1;
    wire stage2_c95_c_fa1;
    wire stage2_c95_s_fa2;
    wire stage2_c95_c_fa2;
    wire stage2_c95_s_fa3;
    wire stage2_c95_c_fa3;
    wire stage2_c96_s_fa0;
    wire stage2_c96_c_fa0;
    wire stage2_c96_s_fa1;
    wire stage2_c96_c_fa1;
    wire stage2_c96_s_fa2;
    wire stage2_c96_c_fa2;
    wire stage2_c96_s_fa3;
    wire stage2_c96_c_fa3;
    wire stage2_c97_s_fa0;
    wire stage2_c97_c_fa0;
    wire stage2_c97_s_fa1;
    wire stage2_c97_c_fa1;
    wire stage2_c97_s_fa2;
    wire stage2_c97_c_fa2;
    wire stage2_c98_s_fa0;
    wire stage2_c98_c_fa0;
    wire stage2_c98_s_fa1;
    wire stage2_c98_c_fa1;
    wire stage2_c98_s_fa2;
    wire stage2_c98_c_fa2;
    wire stage2_c99_s_fa0;
    wire stage2_c99_c_fa0;
    wire stage2_c99_s_fa1;
    wire stage2_c99_c_fa1;
    wire stage2_c99_s_fa2;
    wire stage2_c99_c_fa2;
    wire stage2_c100_s_fa0;
    wire stage2_c100_c_fa0;
    wire stage2_c100_s_fa1;
    wire stage2_c100_c_fa1;
    wire stage2_c100_s_ha0;
    wire stage2_c100_c_ha0;
    wire stage2_c101_s_fa0;
    wire stage2_c101_c_fa0;
    wire stage2_c101_s_fa1;
    wire stage2_c101_c_fa1;
    wire stage2_c101_s_ha0;
    wire stage2_c101_c_ha0;
    wire stage2_c102_s_fa0;
    wire stage2_c102_c_fa0;
    wire stage2_c102_s_fa1;
    wire stage2_c102_c_fa1;
    wire stage2_c102_s_ha0;
    wire stage2_c102_c_ha0;
    wire stage2_c103_s_fa0;
    wire stage2_c103_c_fa0;
    wire stage2_c103_s_fa1;
    wire stage2_c103_c_fa1;
    wire stage2_c104_s_fa0;
    wire stage2_c104_c_fa0;
    wire stage2_c104_s_fa1;
    wire stage2_c104_c_fa1;
    wire stage2_c105_s_fa0;
    wire stage2_c105_c_fa0;
    wire stage2_c105_s_fa1;
    wire stage2_c105_c_fa1;
    wire stage2_c106_s_fa0;
    wire stage2_c106_c_fa0;
    wire stage2_c107_s_fa0;
    wire stage2_c107_c_fa0;
    wire stage2_c108_s_fa0;
    wire stage2_c108_c_fa0;
    wire stage2_c109_s_ha0;
    wire stage2_c109_c_ha0;
    wire stage2_c110_s_ha0;
    wire stage2_c110_c_ha0;
    wire stage2_c111_s_ha0;
    wire stage2_c111_c_ha0;
    wire stage3_c3_s_ha0;
    wire stage3_c3_c_ha0;
    wire stage3_c4_s_ha0;
    wire stage3_c4_c_ha0;
    wire stage3_c5_s_fa0;
    wire stage3_c5_c_fa0;
    wire stage3_c6_s_fa0;
    wire stage3_c6_c_fa0;
    wire stage3_c7_s_fa0;
    wire stage3_c7_c_fa0;
    wire stage3_c8_s_fa0;
    wire stage3_c8_c_fa0;
    wire stage3_c9_s_fa0;
    wire stage3_c9_c_fa0;
    wire stage3_c9_s_ha0;
    wire stage3_c9_c_ha0;
    wire stage3_c10_s_fa0;
    wire stage3_c10_c_fa0;
    wire stage3_c10_s_ha0;
    wire stage3_c10_c_ha0;
    wire stage3_c11_s_fa0;
    wire stage3_c11_c_fa0;
    wire stage3_c11_s_ha0;
    wire stage3_c11_c_ha0;
    wire stage3_c12_s_fa0;
    wire stage3_c12_c_fa0;
    wire stage3_c12_s_fa1;
    wire stage3_c12_c_fa1;
    wire stage3_c13_s_fa0;
    wire stage3_c13_c_fa0;
    wire stage3_c13_s_fa1;
    wire stage3_c13_c_fa1;
    wire stage3_c14_s_fa0;
    wire stage3_c14_c_fa0;
    wire stage3_c14_s_fa1;
    wire stage3_c14_c_fa1;
    wire stage3_c15_s_fa0;
    wire stage3_c15_c_fa0;
    wire stage3_c15_s_fa1;
    wire stage3_c15_c_fa1;
    wire stage3_c16_s_fa0;
    wire stage3_c16_c_fa0;
    wire stage3_c16_s_fa1;
    wire stage3_c16_c_fa1;
    wire stage3_c16_s_ha0;
    wire stage3_c16_c_ha0;
    wire stage3_c17_s_fa0;
    wire stage3_c17_c_fa0;
    wire stage3_c17_s_fa1;
    wire stage3_c17_c_fa1;
    wire stage3_c17_s_ha0;
    wire stage3_c17_c_ha0;
    wire stage3_c18_s_fa0;
    wire stage3_c18_c_fa0;
    wire stage3_c18_s_fa1;
    wire stage3_c18_c_fa1;
    wire stage3_c18_s_fa2;
    wire stage3_c18_c_fa2;
    wire stage3_c19_s_fa0;
    wire stage3_c19_c_fa0;
    wire stage3_c19_s_fa1;
    wire stage3_c19_c_fa1;
    wire stage3_c19_s_fa2;
    wire stage3_c19_c_fa2;
    wire stage3_c20_s_fa0;
    wire stage3_c20_c_fa0;
    wire stage3_c20_s_fa1;
    wire stage3_c20_c_fa1;
    wire stage3_c20_s_fa2;
    wire stage3_c20_c_fa2;
    wire stage3_c21_s_fa0;
    wire stage3_c21_c_fa0;
    wire stage3_c21_s_fa1;
    wire stage3_c21_c_fa1;
    wire stage3_c21_s_fa2;
    wire stage3_c21_c_fa2;
    wire stage3_c22_s_fa0;
    wire stage3_c22_c_fa0;
    wire stage3_c22_s_fa1;
    wire stage3_c22_c_fa1;
    wire stage3_c22_s_fa2;
    wire stage3_c22_c_fa2;
    wire stage3_c23_s_fa0;
    wire stage3_c23_c_fa0;
    wire stage3_c23_s_fa1;
    wire stage3_c23_c_fa1;
    wire stage3_c23_s_fa2;
    wire stage3_c23_c_fa2;
    wire stage3_c23_s_ha0;
    wire stage3_c23_c_ha0;
    wire stage3_c24_s_fa0;
    wire stage3_c24_c_fa0;
    wire stage3_c24_s_fa1;
    wire stage3_c24_c_fa1;
    wire stage3_c24_s_fa2;
    wire stage3_c24_c_fa2;
    wire stage3_c24_s_ha0;
    wire stage3_c24_c_ha0;
    wire stage3_c25_s_fa0;
    wire stage3_c25_c_fa0;
    wire stage3_c25_s_fa1;
    wire stage3_c25_c_fa1;
    wire stage3_c25_s_fa2;
    wire stage3_c25_c_fa2;
    wire stage3_c25_s_fa3;
    wire stage3_c25_c_fa3;
    wire stage3_c26_s_fa0;
    wire stage3_c26_c_fa0;
    wire stage3_c26_s_fa1;
    wire stage3_c26_c_fa1;
    wire stage3_c26_s_fa2;
    wire stage3_c26_c_fa2;
    wire stage3_c26_s_fa3;
    wire stage3_c26_c_fa3;
    wire stage3_c27_s_fa0;
    wire stage3_c27_c_fa0;
    wire stage3_c27_s_fa1;
    wire stage3_c27_c_fa1;
    wire stage3_c27_s_fa2;
    wire stage3_c27_c_fa2;
    wire stage3_c27_s_fa3;
    wire stage3_c27_c_fa3;
    wire stage3_c28_s_fa0;
    wire stage3_c28_c_fa0;
    wire stage3_c28_s_fa1;
    wire stage3_c28_c_fa1;
    wire stage3_c28_s_fa2;
    wire stage3_c28_c_fa2;
    wire stage3_c28_s_fa3;
    wire stage3_c28_c_fa3;
    wire stage3_c29_s_fa0;
    wire stage3_c29_c_fa0;
    wire stage3_c29_s_fa1;
    wire stage3_c29_c_fa1;
    wire stage3_c29_s_fa2;
    wire stage3_c29_c_fa2;
    wire stage3_c29_s_fa3;
    wire stage3_c29_c_fa3;
    wire stage3_c30_s_fa0;
    wire stage3_c30_c_fa0;
    wire stage3_c30_s_fa1;
    wire stage3_c30_c_fa1;
    wire stage3_c30_s_fa2;
    wire stage3_c30_c_fa2;
    wire stage3_c30_s_fa3;
    wire stage3_c30_c_fa3;
    wire stage3_c30_s_ha0;
    wire stage3_c30_c_ha0;
    wire stage3_c31_s_fa0;
    wire stage3_c31_c_fa0;
    wire stage3_c31_s_fa1;
    wire stage3_c31_c_fa1;
    wire stage3_c31_s_fa2;
    wire stage3_c31_c_fa2;
    wire stage3_c31_s_fa3;
    wire stage3_c31_c_fa3;
    wire stage3_c31_s_ha0;
    wire stage3_c31_c_ha0;
    wire stage3_c32_s_fa0;
    wire stage3_c32_c_fa0;
    wire stage3_c32_s_fa1;
    wire stage3_c32_c_fa1;
    wire stage3_c32_s_fa2;
    wire stage3_c32_c_fa2;
    wire stage3_c32_s_fa3;
    wire stage3_c32_c_fa3;
    wire stage3_c32_s_fa4;
    wire stage3_c32_c_fa4;
    wire stage3_c33_s_fa0;
    wire stage3_c33_c_fa0;
    wire stage3_c33_s_fa1;
    wire stage3_c33_c_fa1;
    wire stage3_c33_s_fa2;
    wire stage3_c33_c_fa2;
    wire stage3_c33_s_fa3;
    wire stage3_c33_c_fa3;
    wire stage3_c33_s_fa4;
    wire stage3_c33_c_fa4;
    wire stage3_c34_s_fa0;
    wire stage3_c34_c_fa0;
    wire stage3_c34_s_fa1;
    wire stage3_c34_c_fa1;
    wire stage3_c34_s_fa2;
    wire stage3_c34_c_fa2;
    wire stage3_c34_s_fa3;
    wire stage3_c34_c_fa3;
    wire stage3_c34_s_fa4;
    wire stage3_c34_c_fa4;
    wire stage3_c35_s_fa0;
    wire stage3_c35_c_fa0;
    wire stage3_c35_s_fa1;
    wire stage3_c35_c_fa1;
    wire stage3_c35_s_fa2;
    wire stage3_c35_c_fa2;
    wire stage3_c35_s_fa3;
    wire stage3_c35_c_fa3;
    wire stage3_c35_s_fa4;
    wire stage3_c35_c_fa4;
    wire stage3_c36_s_fa0;
    wire stage3_c36_c_fa0;
    wire stage3_c36_s_fa1;
    wire stage3_c36_c_fa1;
    wire stage3_c36_s_fa2;
    wire stage3_c36_c_fa2;
    wire stage3_c36_s_fa3;
    wire stage3_c36_c_fa3;
    wire stage3_c36_s_fa4;
    wire stage3_c36_c_fa4;
    wire stage3_c36_s_ha0;
    wire stage3_c36_c_ha0;
    wire stage3_c37_s_fa0;
    wire stage3_c37_c_fa0;
    wire stage3_c37_s_fa1;
    wire stage3_c37_c_fa1;
    wire stage3_c37_s_fa2;
    wire stage3_c37_c_fa2;
    wire stage3_c37_s_fa3;
    wire stage3_c37_c_fa3;
    wire stage3_c37_s_fa4;
    wire stage3_c37_c_fa4;
    wire stage3_c37_s_ha0;
    wire stage3_c37_c_ha0;
    wire stage3_c38_s_fa0;
    wire stage3_c38_c_fa0;
    wire stage3_c38_s_fa1;
    wire stage3_c38_c_fa1;
    wire stage3_c38_s_fa2;
    wire stage3_c38_c_fa2;
    wire stage3_c38_s_fa3;
    wire stage3_c38_c_fa3;
    wire stage3_c38_s_fa4;
    wire stage3_c38_c_fa4;
    wire stage3_c38_s_ha0;
    wire stage3_c38_c_ha0;
    wire stage3_c39_s_fa0;
    wire stage3_c39_c_fa0;
    wire stage3_c39_s_fa1;
    wire stage3_c39_c_fa1;
    wire stage3_c39_s_fa2;
    wire stage3_c39_c_fa2;
    wire stage3_c39_s_fa3;
    wire stage3_c39_c_fa3;
    wire stage3_c39_s_fa4;
    wire stage3_c39_c_fa4;
    wire stage3_c39_s_fa5;
    wire stage3_c39_c_fa5;
    wire stage3_c40_s_fa0;
    wire stage3_c40_c_fa0;
    wire stage3_c40_s_fa1;
    wire stage3_c40_c_fa1;
    wire stage3_c40_s_fa2;
    wire stage3_c40_c_fa2;
    wire stage3_c40_s_fa3;
    wire stage3_c40_c_fa3;
    wire stage3_c40_s_fa4;
    wire stage3_c40_c_fa4;
    wire stage3_c40_s_fa5;
    wire stage3_c40_c_fa5;
    wire stage3_c41_s_fa0;
    wire stage3_c41_c_fa0;
    wire stage3_c41_s_fa1;
    wire stage3_c41_c_fa1;
    wire stage3_c41_s_fa2;
    wire stage3_c41_c_fa2;
    wire stage3_c41_s_fa3;
    wire stage3_c41_c_fa3;
    wire stage3_c41_s_fa4;
    wire stage3_c41_c_fa4;
    wire stage3_c41_s_fa5;
    wire stage3_c41_c_fa5;
    wire stage3_c42_s_fa0;
    wire stage3_c42_c_fa0;
    wire stage3_c42_s_fa1;
    wire stage3_c42_c_fa1;
    wire stage3_c42_s_fa2;
    wire stage3_c42_c_fa2;
    wire stage3_c42_s_fa3;
    wire stage3_c42_c_fa3;
    wire stage3_c42_s_fa4;
    wire stage3_c42_c_fa4;
    wire stage3_c42_s_fa5;
    wire stage3_c42_c_fa5;
    wire stage3_c43_s_fa0;
    wire stage3_c43_c_fa0;
    wire stage3_c43_s_fa1;
    wire stage3_c43_c_fa1;
    wire stage3_c43_s_fa2;
    wire stage3_c43_c_fa2;
    wire stage3_c43_s_fa3;
    wire stage3_c43_c_fa3;
    wire stage3_c43_s_fa4;
    wire stage3_c43_c_fa4;
    wire stage3_c43_s_fa5;
    wire stage3_c43_c_fa5;
    wire stage3_c44_s_fa0;
    wire stage3_c44_c_fa0;
    wire stage3_c44_s_fa1;
    wire stage3_c44_c_fa1;
    wire stage3_c44_s_fa2;
    wire stage3_c44_c_fa2;
    wire stage3_c44_s_fa3;
    wire stage3_c44_c_fa3;
    wire stage3_c44_s_fa4;
    wire stage3_c44_c_fa4;
    wire stage3_c44_s_fa5;
    wire stage3_c44_c_fa5;
    wire stage3_c45_s_fa0;
    wire stage3_c45_c_fa0;
    wire stage3_c45_s_fa1;
    wire stage3_c45_c_fa1;
    wire stage3_c45_s_fa2;
    wire stage3_c45_c_fa2;
    wire stage3_c45_s_fa3;
    wire stage3_c45_c_fa3;
    wire stage3_c45_s_fa4;
    wire stage3_c45_c_fa4;
    wire stage3_c45_s_fa5;
    wire stage3_c45_c_fa5;
    wire stage3_c46_s_fa0;
    wire stage3_c46_c_fa0;
    wire stage3_c46_s_fa1;
    wire stage3_c46_c_fa1;
    wire stage3_c46_s_fa2;
    wire stage3_c46_c_fa2;
    wire stage3_c46_s_fa3;
    wire stage3_c46_c_fa3;
    wire stage3_c46_s_fa4;
    wire stage3_c46_c_fa4;
    wire stage3_c46_s_fa5;
    wire stage3_c46_c_fa5;
    wire stage3_c47_s_fa0;
    wire stage3_c47_c_fa0;
    wire stage3_c47_s_fa1;
    wire stage3_c47_c_fa1;
    wire stage3_c47_s_fa2;
    wire stage3_c47_c_fa2;
    wire stage3_c47_s_fa3;
    wire stage3_c47_c_fa3;
    wire stage3_c47_s_fa4;
    wire stage3_c47_c_fa4;
    wire stage3_c47_s_fa5;
    wire stage3_c47_c_fa5;
    wire stage3_c48_s_fa0;
    wire stage3_c48_c_fa0;
    wire stage3_c48_s_fa1;
    wire stage3_c48_c_fa1;
    wire stage3_c48_s_fa2;
    wire stage3_c48_c_fa2;
    wire stage3_c48_s_fa3;
    wire stage3_c48_c_fa3;
    wire stage3_c48_s_fa4;
    wire stage3_c48_c_fa4;
    wire stage3_c48_s_fa5;
    wire stage3_c48_c_fa5;
    wire stage3_c49_s_fa0;
    wire stage3_c49_c_fa0;
    wire stage3_c49_s_fa1;
    wire stage3_c49_c_fa1;
    wire stage3_c49_s_fa2;
    wire stage3_c49_c_fa2;
    wire stage3_c49_s_fa3;
    wire stage3_c49_c_fa3;
    wire stage3_c49_s_fa4;
    wire stage3_c49_c_fa4;
    wire stage3_c49_s_fa5;
    wire stage3_c49_c_fa5;
    wire stage3_c50_s_fa0;
    wire stage3_c50_c_fa0;
    wire stage3_c50_s_fa1;
    wire stage3_c50_c_fa1;
    wire stage3_c50_s_fa2;
    wire stage3_c50_c_fa2;
    wire stage3_c50_s_fa3;
    wire stage3_c50_c_fa3;
    wire stage3_c50_s_fa4;
    wire stage3_c50_c_fa4;
    wire stage3_c50_s_fa5;
    wire stage3_c50_c_fa5;
    wire stage3_c51_s_fa0;
    wire stage3_c51_c_fa0;
    wire stage3_c51_s_fa1;
    wire stage3_c51_c_fa1;
    wire stage3_c51_s_fa2;
    wire stage3_c51_c_fa2;
    wire stage3_c51_s_fa3;
    wire stage3_c51_c_fa3;
    wire stage3_c51_s_fa4;
    wire stage3_c51_c_fa4;
    wire stage3_c51_s_fa5;
    wire stage3_c51_c_fa5;
    wire stage3_c52_s_fa0;
    wire stage3_c52_c_fa0;
    wire stage3_c52_s_fa1;
    wire stage3_c52_c_fa1;
    wire stage3_c52_s_fa2;
    wire stage3_c52_c_fa2;
    wire stage3_c52_s_fa3;
    wire stage3_c52_c_fa3;
    wire stage3_c52_s_fa4;
    wire stage3_c52_c_fa4;
    wire stage3_c52_s_fa5;
    wire stage3_c52_c_fa5;
    wire stage3_c53_s_fa0;
    wire stage3_c53_c_fa0;
    wire stage3_c53_s_fa1;
    wire stage3_c53_c_fa1;
    wire stage3_c53_s_fa2;
    wire stage3_c53_c_fa2;
    wire stage3_c53_s_fa3;
    wire stage3_c53_c_fa3;
    wire stage3_c53_s_fa4;
    wire stage3_c53_c_fa4;
    wire stage3_c53_s_fa5;
    wire stage3_c53_c_fa5;
    wire stage3_c54_s_fa0;
    wire stage3_c54_c_fa0;
    wire stage3_c54_s_fa1;
    wire stage3_c54_c_fa1;
    wire stage3_c54_s_fa2;
    wire stage3_c54_c_fa2;
    wire stage3_c54_s_fa3;
    wire stage3_c54_c_fa3;
    wire stage3_c54_s_fa4;
    wire stage3_c54_c_fa4;
    wire stage3_c54_s_fa5;
    wire stage3_c54_c_fa5;
    wire stage3_c55_s_fa0;
    wire stage3_c55_c_fa0;
    wire stage3_c55_s_fa1;
    wire stage3_c55_c_fa1;
    wire stage3_c55_s_fa2;
    wire stage3_c55_c_fa2;
    wire stage3_c55_s_fa3;
    wire stage3_c55_c_fa3;
    wire stage3_c55_s_fa4;
    wire stage3_c55_c_fa4;
    wire stage3_c55_s_fa5;
    wire stage3_c55_c_fa5;
    wire stage3_c56_s_fa0;
    wire stage3_c56_c_fa0;
    wire stage3_c56_s_fa1;
    wire stage3_c56_c_fa1;
    wire stage3_c56_s_fa2;
    wire stage3_c56_c_fa2;
    wire stage3_c56_s_fa3;
    wire stage3_c56_c_fa3;
    wire stage3_c56_s_fa4;
    wire stage3_c56_c_fa4;
    wire stage3_c56_s_fa5;
    wire stage3_c56_c_fa5;
    wire stage3_c57_s_fa0;
    wire stage3_c57_c_fa0;
    wire stage3_c57_s_fa1;
    wire stage3_c57_c_fa1;
    wire stage3_c57_s_fa2;
    wire stage3_c57_c_fa2;
    wire stage3_c57_s_fa3;
    wire stage3_c57_c_fa3;
    wire stage3_c57_s_fa4;
    wire stage3_c57_c_fa4;
    wire stage3_c57_s_fa5;
    wire stage3_c57_c_fa5;
    wire stage3_c58_s_fa0;
    wire stage3_c58_c_fa0;
    wire stage3_c58_s_fa1;
    wire stage3_c58_c_fa1;
    wire stage3_c58_s_fa2;
    wire stage3_c58_c_fa2;
    wire stage3_c58_s_fa3;
    wire stage3_c58_c_fa3;
    wire stage3_c58_s_fa4;
    wire stage3_c58_c_fa4;
    wire stage3_c58_s_fa5;
    wire stage3_c58_c_fa5;
    wire stage3_c59_s_fa0;
    wire stage3_c59_c_fa0;
    wire stage3_c59_s_fa1;
    wire stage3_c59_c_fa1;
    wire stage3_c59_s_fa2;
    wire stage3_c59_c_fa2;
    wire stage3_c59_s_fa3;
    wire stage3_c59_c_fa3;
    wire stage3_c59_s_fa4;
    wire stage3_c59_c_fa4;
    wire stage3_c59_s_fa5;
    wire stage3_c59_c_fa5;
    wire stage3_c60_s_fa0;
    wire stage3_c60_c_fa0;
    wire stage3_c60_s_fa1;
    wire stage3_c60_c_fa1;
    wire stage3_c60_s_fa2;
    wire stage3_c60_c_fa2;
    wire stage3_c60_s_fa3;
    wire stage3_c60_c_fa3;
    wire stage3_c60_s_fa4;
    wire stage3_c60_c_fa4;
    wire stage3_c60_s_fa5;
    wire stage3_c60_c_fa5;
    wire stage3_c61_s_fa0;
    wire stage3_c61_c_fa0;
    wire stage3_c61_s_fa1;
    wire stage3_c61_c_fa1;
    wire stage3_c61_s_fa2;
    wire stage3_c61_c_fa2;
    wire stage3_c61_s_fa3;
    wire stage3_c61_c_fa3;
    wire stage3_c61_s_fa4;
    wire stage3_c61_c_fa4;
    wire stage3_c61_s_fa5;
    wire stage3_c61_c_fa5;
    wire stage3_c62_s_fa0;
    wire stage3_c62_c_fa0;
    wire stage3_c62_s_fa1;
    wire stage3_c62_c_fa1;
    wire stage3_c62_s_fa2;
    wire stage3_c62_c_fa2;
    wire stage3_c62_s_fa3;
    wire stage3_c62_c_fa3;
    wire stage3_c62_s_fa4;
    wire stage3_c62_c_fa4;
    wire stage3_c62_s_fa5;
    wire stage3_c62_c_fa5;
    wire stage3_c63_s_fa0;
    wire stage3_c63_c_fa0;
    wire stage3_c63_s_fa1;
    wire stage3_c63_c_fa1;
    wire stage3_c63_s_fa2;
    wire stage3_c63_c_fa2;
    wire stage3_c63_s_fa3;
    wire stage3_c63_c_fa3;
    wire stage3_c63_s_fa4;
    wire stage3_c63_c_fa4;
    wire stage3_c63_s_fa5;
    wire stage3_c63_c_fa5;
    wire stage3_c64_s_fa0;
    wire stage3_c64_c_fa0;
    wire stage3_c64_s_fa1;
    wire stage3_c64_c_fa1;
    wire stage3_c64_s_fa2;
    wire stage3_c64_c_fa2;
    wire stage3_c64_s_fa3;
    wire stage3_c64_c_fa3;
    wire stage3_c64_s_fa4;
    wire stage3_c64_c_fa4;
    wire stage3_c64_s_fa5;
    wire stage3_c64_c_fa5;
    wire stage3_c65_s_fa0;
    wire stage3_c65_c_fa0;
    wire stage3_c65_s_fa1;
    wire stage3_c65_c_fa1;
    wire stage3_c65_s_fa2;
    wire stage3_c65_c_fa2;
    wire stage3_c65_s_fa3;
    wire stage3_c65_c_fa3;
    wire stage3_c65_s_fa4;
    wire stage3_c65_c_fa4;
    wire stage3_c65_s_fa5;
    wire stage3_c65_c_fa5;
    wire stage3_c66_s_fa0;
    wire stage3_c66_c_fa0;
    wire stage3_c66_s_fa1;
    wire stage3_c66_c_fa1;
    wire stage3_c66_s_fa2;
    wire stage3_c66_c_fa2;
    wire stage3_c66_s_fa3;
    wire stage3_c66_c_fa3;
    wire stage3_c66_s_fa4;
    wire stage3_c66_c_fa4;
    wire stage3_c66_s_fa5;
    wire stage3_c66_c_fa5;
    wire stage3_c67_s_fa0;
    wire stage3_c67_c_fa0;
    wire stage3_c67_s_fa1;
    wire stage3_c67_c_fa1;
    wire stage3_c67_s_fa2;
    wire stage3_c67_c_fa2;
    wire stage3_c67_s_fa3;
    wire stage3_c67_c_fa3;
    wire stage3_c67_s_fa4;
    wire stage3_c67_c_fa4;
    wire stage3_c67_s_fa5;
    wire stage3_c67_c_fa5;
    wire stage3_c68_s_fa0;
    wire stage3_c68_c_fa0;
    wire stage3_c68_s_fa1;
    wire stage3_c68_c_fa1;
    wire stage3_c68_s_fa2;
    wire stage3_c68_c_fa2;
    wire stage3_c68_s_fa3;
    wire stage3_c68_c_fa3;
    wire stage3_c68_s_fa4;
    wire stage3_c68_c_fa4;
    wire stage3_c68_s_fa5;
    wire stage3_c68_c_fa5;
    wire stage3_c69_s_fa0;
    wire stage3_c69_c_fa0;
    wire stage3_c69_s_fa1;
    wire stage3_c69_c_fa1;
    wire stage3_c69_s_fa2;
    wire stage3_c69_c_fa2;
    wire stage3_c69_s_fa3;
    wire stage3_c69_c_fa3;
    wire stage3_c69_s_fa4;
    wire stage3_c69_c_fa4;
    wire stage3_c69_s_fa5;
    wire stage3_c69_c_fa5;
    wire stage3_c70_s_fa0;
    wire stage3_c70_c_fa0;
    wire stage3_c70_s_fa1;
    wire stage3_c70_c_fa1;
    wire stage3_c70_s_fa2;
    wire stage3_c70_c_fa2;
    wire stage3_c70_s_fa3;
    wire stage3_c70_c_fa3;
    wire stage3_c70_s_fa4;
    wire stage3_c70_c_fa4;
    wire stage3_c70_s_fa5;
    wire stage3_c70_c_fa5;
    wire stage3_c71_s_fa0;
    wire stage3_c71_c_fa0;
    wire stage3_c71_s_fa1;
    wire stage3_c71_c_fa1;
    wire stage3_c71_s_fa2;
    wire stage3_c71_c_fa2;
    wire stage3_c71_s_fa3;
    wire stage3_c71_c_fa3;
    wire stage3_c71_s_fa4;
    wire stage3_c71_c_fa4;
    wire stage3_c71_s_fa5;
    wire stage3_c71_c_fa5;
    wire stage3_c72_s_fa0;
    wire stage3_c72_c_fa0;
    wire stage3_c72_s_fa1;
    wire stage3_c72_c_fa1;
    wire stage3_c72_s_fa2;
    wire stage3_c72_c_fa2;
    wire stage3_c72_s_fa3;
    wire stage3_c72_c_fa3;
    wire stage3_c72_s_fa4;
    wire stage3_c72_c_fa4;
    wire stage3_c72_s_fa5;
    wire stage3_c72_c_fa5;
    wire stage3_c73_s_fa0;
    wire stage3_c73_c_fa0;
    wire stage3_c73_s_fa1;
    wire stage3_c73_c_fa1;
    wire stage3_c73_s_fa2;
    wire stage3_c73_c_fa2;
    wire stage3_c73_s_fa3;
    wire stage3_c73_c_fa3;
    wire stage3_c73_s_fa4;
    wire stage3_c73_c_fa4;
    wire stage3_c73_s_fa5;
    wire stage3_c73_c_fa5;
    wire stage3_c74_s_fa0;
    wire stage3_c74_c_fa0;
    wire stage3_c74_s_fa1;
    wire stage3_c74_c_fa1;
    wire stage3_c74_s_fa2;
    wire stage3_c74_c_fa2;
    wire stage3_c74_s_fa3;
    wire stage3_c74_c_fa3;
    wire stage3_c74_s_fa4;
    wire stage3_c74_c_fa4;
    wire stage3_c74_s_fa5;
    wire stage3_c74_c_fa5;
    wire stage3_c75_s_fa0;
    wire stage3_c75_c_fa0;
    wire stage3_c75_s_fa1;
    wire stage3_c75_c_fa1;
    wire stage3_c75_s_fa2;
    wire stage3_c75_c_fa2;
    wire stage3_c75_s_fa3;
    wire stage3_c75_c_fa3;
    wire stage3_c75_s_fa4;
    wire stage3_c75_c_fa4;
    wire stage3_c75_s_fa5;
    wire stage3_c75_c_fa5;
    wire stage3_c76_s_fa0;
    wire stage3_c76_c_fa0;
    wire stage3_c76_s_fa1;
    wire stage3_c76_c_fa1;
    wire stage3_c76_s_fa2;
    wire stage3_c76_c_fa2;
    wire stage3_c76_s_fa3;
    wire stage3_c76_c_fa3;
    wire stage3_c76_s_fa4;
    wire stage3_c76_c_fa4;
    wire stage3_c76_s_ha0;
    wire stage3_c76_c_ha0;
    wire stage3_c77_s_fa0;
    wire stage3_c77_c_fa0;
    wire stage3_c77_s_fa1;
    wire stage3_c77_c_fa1;
    wire stage3_c77_s_fa2;
    wire stage3_c77_c_fa2;
    wire stage3_c77_s_fa3;
    wire stage3_c77_c_fa3;
    wire stage3_c77_s_fa4;
    wire stage3_c77_c_fa4;
    wire stage3_c78_s_fa0;
    wire stage3_c78_c_fa0;
    wire stage3_c78_s_fa1;
    wire stage3_c78_c_fa1;
    wire stage3_c78_s_fa2;
    wire stage3_c78_c_fa2;
    wire stage3_c78_s_fa3;
    wire stage3_c78_c_fa3;
    wire stage3_c78_s_fa4;
    wire stage3_c78_c_fa4;
    wire stage3_c79_s_fa0;
    wire stage3_c79_c_fa0;
    wire stage3_c79_s_fa1;
    wire stage3_c79_c_fa1;
    wire stage3_c79_s_fa2;
    wire stage3_c79_c_fa2;
    wire stage3_c79_s_fa3;
    wire stage3_c79_c_fa3;
    wire stage3_c79_s_fa4;
    wire stage3_c79_c_fa4;
    wire stage3_c80_s_fa0;
    wire stage3_c80_c_fa0;
    wire stage3_c80_s_fa1;
    wire stage3_c80_c_fa1;
    wire stage3_c80_s_fa2;
    wire stage3_c80_c_fa2;
    wire stage3_c80_s_fa3;
    wire stage3_c80_c_fa3;
    wire stage3_c80_s_fa4;
    wire stage3_c80_c_fa4;
    wire stage3_c81_s_fa0;
    wire stage3_c81_c_fa0;
    wire stage3_c81_s_fa1;
    wire stage3_c81_c_fa1;
    wire stage3_c81_s_fa2;
    wire stage3_c81_c_fa2;
    wire stage3_c81_s_fa3;
    wire stage3_c81_c_fa3;
    wire stage3_c81_s_fa4;
    wire stage3_c81_c_fa4;
    wire stage3_c82_s_fa0;
    wire stage3_c82_c_fa0;
    wire stage3_c82_s_fa1;
    wire stage3_c82_c_fa1;
    wire stage3_c82_s_fa2;
    wire stage3_c82_c_fa2;
    wire stage3_c82_s_fa3;
    wire stage3_c82_c_fa3;
    wire stage3_c82_s_ha0;
    wire stage3_c82_c_ha0;
    wire stage3_c83_s_fa0;
    wire stage3_c83_c_fa0;
    wire stage3_c83_s_fa1;
    wire stage3_c83_c_fa1;
    wire stage3_c83_s_fa2;
    wire stage3_c83_c_fa2;
    wire stage3_c83_s_fa3;
    wire stage3_c83_c_fa3;
    wire stage3_c83_s_ha0;
    wire stage3_c83_c_ha0;
    wire stage3_c84_s_fa0;
    wire stage3_c84_c_fa0;
    wire stage3_c84_s_fa1;
    wire stage3_c84_c_fa1;
    wire stage3_c84_s_fa2;
    wire stage3_c84_c_fa2;
    wire stage3_c84_s_fa3;
    wire stage3_c84_c_fa3;
    wire stage3_c84_s_ha0;
    wire stage3_c84_c_ha0;
    wire stage3_c85_s_fa0;
    wire stage3_c85_c_fa0;
    wire stage3_c85_s_fa1;
    wire stage3_c85_c_fa1;
    wire stage3_c85_s_fa2;
    wire stage3_c85_c_fa2;
    wire stage3_c85_s_fa3;
    wire stage3_c85_c_fa3;
    wire stage3_c86_s_fa0;
    wire stage3_c86_c_fa0;
    wire stage3_c86_s_fa1;
    wire stage3_c86_c_fa1;
    wire stage3_c86_s_fa2;
    wire stage3_c86_c_fa2;
    wire stage3_c86_s_fa3;
    wire stage3_c86_c_fa3;
    wire stage3_c87_s_fa0;
    wire stage3_c87_c_fa0;
    wire stage3_c87_s_fa1;
    wire stage3_c87_c_fa1;
    wire stage3_c87_s_fa2;
    wire stage3_c87_c_fa2;
    wire stage3_c87_s_fa3;
    wire stage3_c87_c_fa3;
    wire stage3_c88_s_fa0;
    wire stage3_c88_c_fa0;
    wire stage3_c88_s_fa1;
    wire stage3_c88_c_fa1;
    wire stage3_c88_s_fa2;
    wire stage3_c88_c_fa2;
    wire stage3_c88_s_fa3;
    wire stage3_c88_c_fa3;
    wire stage3_c89_s_fa0;
    wire stage3_c89_c_fa0;
    wire stage3_c89_s_fa1;
    wire stage3_c89_c_fa1;
    wire stage3_c89_s_fa2;
    wire stage3_c89_c_fa2;
    wire stage3_c89_s_ha0;
    wire stage3_c89_c_ha0;
    wire stage3_c90_s_fa0;
    wire stage3_c90_c_fa0;
    wire stage3_c90_s_fa1;
    wire stage3_c90_c_fa1;
    wire stage3_c90_s_fa2;
    wire stage3_c90_c_fa2;
    wire stage3_c90_s_ha0;
    wire stage3_c90_c_ha0;
    wire stage3_c91_s_fa0;
    wire stage3_c91_c_fa0;
    wire stage3_c91_s_fa1;
    wire stage3_c91_c_fa1;
    wire stage3_c91_s_fa2;
    wire stage3_c91_c_fa2;
    wire stage3_c92_s_fa0;
    wire stage3_c92_c_fa0;
    wire stage3_c92_s_fa1;
    wire stage3_c92_c_fa1;
    wire stage3_c92_s_fa2;
    wire stage3_c92_c_fa2;
    wire stage3_c93_s_fa0;
    wire stage3_c93_c_fa0;
    wire stage3_c93_s_fa1;
    wire stage3_c93_c_fa1;
    wire stage3_c93_s_fa2;
    wire stage3_c93_c_fa2;
    wire stage3_c94_s_fa0;
    wire stage3_c94_c_fa0;
    wire stage3_c94_s_fa1;
    wire stage3_c94_c_fa1;
    wire stage3_c94_s_fa2;
    wire stage3_c94_c_fa2;
    wire stage3_c95_s_fa0;
    wire stage3_c95_c_fa0;
    wire stage3_c95_s_fa1;
    wire stage3_c95_c_fa1;
    wire stage3_c95_s_ha0;
    wire stage3_c95_c_ha0;
    wire stage3_c96_s_fa0;
    wire stage3_c96_c_fa0;
    wire stage3_c96_s_fa1;
    wire stage3_c96_c_fa1;
    wire stage3_c96_s_ha0;
    wire stage3_c96_c_ha0;
    wire stage3_c97_s_fa0;
    wire stage3_c97_c_fa0;
    wire stage3_c97_s_fa1;
    wire stage3_c97_c_fa1;
    wire stage3_c97_s_ha0;
    wire stage3_c97_c_ha0;
    wire stage3_c98_s_fa0;
    wire stage3_c98_c_fa0;
    wire stage3_c98_s_fa1;
    wire stage3_c98_c_fa1;
    wire stage3_c99_s_fa0;
    wire stage3_c99_c_fa0;
    wire stage3_c99_s_fa1;
    wire stage3_c99_c_fa1;
    wire stage3_c100_s_fa0;
    wire stage3_c100_c_fa0;
    wire stage3_c100_s_fa1;
    wire stage3_c100_c_fa1;
    wire stage3_c101_s_fa0;
    wire stage3_c101_c_fa0;
    wire stage3_c101_s_fa1;
    wire stage3_c101_c_fa1;
    wire stage3_c102_s_fa0;
    wire stage3_c102_c_fa0;
    wire stage3_c102_s_fa1;
    wire stage3_c102_c_fa1;
    wire stage3_c103_s_fa0;
    wire stage3_c103_c_fa0;
    wire stage3_c103_s_ha0;
    wire stage3_c103_c_ha0;
    wire stage3_c104_s_fa0;
    wire stage3_c104_c_fa0;
    wire stage3_c105_s_fa0;
    wire stage3_c105_c_fa0;
    wire stage3_c106_s_fa0;
    wire stage3_c106_c_fa0;
    wire stage3_c107_s_fa0;
    wire stage3_c107_c_fa0;
    wire stage3_c108_s_fa0;
    wire stage3_c108_c_fa0;
    wire stage3_c109_s_ha0;
    wire stage3_c109_c_ha0;
    wire stage3_c110_s_ha0;
    wire stage3_c110_c_ha0;
    wire stage3_c111_s_ha0;
    wire stage3_c111_c_ha0;
    wire stage4_c4_s_ha0;
    wire stage4_c4_c_ha0;
    wire stage4_c5_s_ha0;
    wire stage4_c5_c_ha0;
    wire stage4_c6_s_ha0;
    wire stage4_c6_c_ha0;
    wire stage4_c7_s_fa0;
    wire stage4_c7_c_fa0;
    wire stage4_c8_s_fa0;
    wire stage4_c8_c_fa0;
    wire stage4_c9_s_fa0;
    wire stage4_c9_c_fa0;
    wire stage4_c10_s_fa0;
    wire stage4_c10_c_fa0;
    wire stage4_c11_s_fa0;
    wire stage4_c11_c_fa0;
    wire stage4_c12_s_fa0;
    wire stage4_c12_c_fa0;
    wire stage4_c13_s_fa0;
    wire stage4_c13_c_fa0;
    wire stage4_c14_s_fa0;
    wire stage4_c14_c_fa0;
    wire stage4_c14_s_ha0;
    wire stage4_c14_c_ha0;
    wire stage4_c15_s_fa0;
    wire stage4_c15_c_fa0;
    wire stage4_c15_s_ha0;
    wire stage4_c15_c_ha0;
    wire stage4_c16_s_fa0;
    wire stage4_c16_c_fa0;
    wire stage4_c16_s_ha0;
    wire stage4_c16_c_ha0;
    wire stage4_c17_s_fa0;
    wire stage4_c17_c_fa0;
    wire stage4_c17_s_fa1;
    wire stage4_c17_c_fa1;
    wire stage4_c18_s_fa0;
    wire stage4_c18_c_fa0;
    wire stage4_c18_s_fa1;
    wire stage4_c18_c_fa1;
    wire stage4_c19_s_fa0;
    wire stage4_c19_c_fa0;
    wire stage4_c19_s_fa1;
    wire stage4_c19_c_fa1;
    wire stage4_c20_s_fa0;
    wire stage4_c20_c_fa0;
    wire stage4_c20_s_fa1;
    wire stage4_c20_c_fa1;
    wire stage4_c21_s_fa0;
    wire stage4_c21_c_fa0;
    wire stage4_c21_s_fa1;
    wire stage4_c21_c_fa1;
    wire stage4_c22_s_fa0;
    wire stage4_c22_c_fa0;
    wire stage4_c22_s_fa1;
    wire stage4_c22_c_fa1;
    wire stage4_c23_s_fa0;
    wire stage4_c23_c_fa0;
    wire stage4_c23_s_fa1;
    wire stage4_c23_c_fa1;
    wire stage4_c24_s_fa0;
    wire stage4_c24_c_fa0;
    wire stage4_c24_s_fa1;
    wire stage4_c24_c_fa1;
    wire stage4_c24_s_ha0;
    wire stage4_c24_c_ha0;
    wire stage4_c25_s_fa0;
    wire stage4_c25_c_fa0;
    wire stage4_c25_s_fa1;
    wire stage4_c25_c_fa1;
    wire stage4_c25_s_ha0;
    wire stage4_c25_c_ha0;
    wire stage4_c26_s_fa0;
    wire stage4_c26_c_fa0;
    wire stage4_c26_s_fa1;
    wire stage4_c26_c_fa1;
    wire stage4_c26_s_ha0;
    wire stage4_c26_c_ha0;
    wire stage4_c27_s_fa0;
    wire stage4_c27_c_fa0;
    wire stage4_c27_s_fa1;
    wire stage4_c27_c_fa1;
    wire stage4_c27_s_fa2;
    wire stage4_c27_c_fa2;
    wire stage4_c28_s_fa0;
    wire stage4_c28_c_fa0;
    wire stage4_c28_s_fa1;
    wire stage4_c28_c_fa1;
    wire stage4_c28_s_fa2;
    wire stage4_c28_c_fa2;
    wire stage4_c29_s_fa0;
    wire stage4_c29_c_fa0;
    wire stage4_c29_s_fa1;
    wire stage4_c29_c_fa1;
    wire stage4_c29_s_fa2;
    wire stage4_c29_c_fa2;
    wire stage4_c30_s_fa0;
    wire stage4_c30_c_fa0;
    wire stage4_c30_s_fa1;
    wire stage4_c30_c_fa1;
    wire stage4_c30_s_fa2;
    wire stage4_c30_c_fa2;
    wire stage4_c31_s_fa0;
    wire stage4_c31_c_fa0;
    wire stage4_c31_s_fa1;
    wire stage4_c31_c_fa1;
    wire stage4_c31_s_fa2;
    wire stage4_c31_c_fa2;
    wire stage4_c32_s_fa0;
    wire stage4_c32_c_fa0;
    wire stage4_c32_s_fa1;
    wire stage4_c32_c_fa1;
    wire stage4_c32_s_fa2;
    wire stage4_c32_c_fa2;
    wire stage4_c33_s_fa0;
    wire stage4_c33_c_fa0;
    wire stage4_c33_s_fa1;
    wire stage4_c33_c_fa1;
    wire stage4_c33_s_fa2;
    wire stage4_c33_c_fa2;
    wire stage4_c34_s_fa0;
    wire stage4_c34_c_fa0;
    wire stage4_c34_s_fa1;
    wire stage4_c34_c_fa1;
    wire stage4_c34_s_fa2;
    wire stage4_c34_c_fa2;
    wire stage4_c34_s_ha0;
    wire stage4_c34_c_ha0;
    wire stage4_c35_s_fa0;
    wire stage4_c35_c_fa0;
    wire stage4_c35_s_fa1;
    wire stage4_c35_c_fa1;
    wire stage4_c35_s_fa2;
    wire stage4_c35_c_fa2;
    wire stage4_c35_s_ha0;
    wire stage4_c35_c_ha0;
    wire stage4_c36_s_fa0;
    wire stage4_c36_c_fa0;
    wire stage4_c36_s_fa1;
    wire stage4_c36_c_fa1;
    wire stage4_c36_s_fa2;
    wire stage4_c36_c_fa2;
    wire stage4_c36_s_ha0;
    wire stage4_c36_c_ha0;
    wire stage4_c37_s_fa0;
    wire stage4_c37_c_fa0;
    wire stage4_c37_s_fa1;
    wire stage4_c37_c_fa1;
    wire stage4_c37_s_fa2;
    wire stage4_c37_c_fa2;
    wire stage4_c37_s_fa3;
    wire stage4_c37_c_fa3;
    wire stage4_c38_s_fa0;
    wire stage4_c38_c_fa0;
    wire stage4_c38_s_fa1;
    wire stage4_c38_c_fa1;
    wire stage4_c38_s_fa2;
    wire stage4_c38_c_fa2;
    wire stage4_c38_s_fa3;
    wire stage4_c38_c_fa3;
    wire stage4_c39_s_fa0;
    wire stage4_c39_c_fa0;
    wire stage4_c39_s_fa1;
    wire stage4_c39_c_fa1;
    wire stage4_c39_s_fa2;
    wire stage4_c39_c_fa2;
    wire stage4_c39_s_fa3;
    wire stage4_c39_c_fa3;
    wire stage4_c40_s_fa0;
    wire stage4_c40_c_fa0;
    wire stage4_c40_s_fa1;
    wire stage4_c40_c_fa1;
    wire stage4_c40_s_fa2;
    wire stage4_c40_c_fa2;
    wire stage4_c40_s_fa3;
    wire stage4_c40_c_fa3;
    wire stage4_c41_s_fa0;
    wire stage4_c41_c_fa0;
    wire stage4_c41_s_fa1;
    wire stage4_c41_c_fa1;
    wire stage4_c41_s_fa2;
    wire stage4_c41_c_fa2;
    wire stage4_c41_s_fa3;
    wire stage4_c41_c_fa3;
    wire stage4_c42_s_fa0;
    wire stage4_c42_c_fa0;
    wire stage4_c42_s_fa1;
    wire stage4_c42_c_fa1;
    wire stage4_c42_s_fa2;
    wire stage4_c42_c_fa2;
    wire stage4_c42_s_fa3;
    wire stage4_c42_c_fa3;
    wire stage4_c43_s_fa0;
    wire stage4_c43_c_fa0;
    wire stage4_c43_s_fa1;
    wire stage4_c43_c_fa1;
    wire stage4_c43_s_fa2;
    wire stage4_c43_c_fa2;
    wire stage4_c43_s_fa3;
    wire stage4_c43_c_fa3;
    wire stage4_c44_s_fa0;
    wire stage4_c44_c_fa0;
    wire stage4_c44_s_fa1;
    wire stage4_c44_c_fa1;
    wire stage4_c44_s_fa2;
    wire stage4_c44_c_fa2;
    wire stage4_c44_s_fa3;
    wire stage4_c44_c_fa3;
    wire stage4_c45_s_fa0;
    wire stage4_c45_c_fa0;
    wire stage4_c45_s_fa1;
    wire stage4_c45_c_fa1;
    wire stage4_c45_s_fa2;
    wire stage4_c45_c_fa2;
    wire stage4_c45_s_fa3;
    wire stage4_c45_c_fa3;
    wire stage4_c46_s_fa0;
    wire stage4_c46_c_fa0;
    wire stage4_c46_s_fa1;
    wire stage4_c46_c_fa1;
    wire stage4_c46_s_fa2;
    wire stage4_c46_c_fa2;
    wire stage4_c46_s_fa3;
    wire stage4_c46_c_fa3;
    wire stage4_c47_s_fa0;
    wire stage4_c47_c_fa0;
    wire stage4_c47_s_fa1;
    wire stage4_c47_c_fa1;
    wire stage4_c47_s_fa2;
    wire stage4_c47_c_fa2;
    wire stage4_c47_s_fa3;
    wire stage4_c47_c_fa3;
    wire stage4_c48_s_fa0;
    wire stage4_c48_c_fa0;
    wire stage4_c48_s_fa1;
    wire stage4_c48_c_fa1;
    wire stage4_c48_s_fa2;
    wire stage4_c48_c_fa2;
    wire stage4_c48_s_fa3;
    wire stage4_c48_c_fa3;
    wire stage4_c49_s_fa0;
    wire stage4_c49_c_fa0;
    wire stage4_c49_s_fa1;
    wire stage4_c49_c_fa1;
    wire stage4_c49_s_fa2;
    wire stage4_c49_c_fa2;
    wire stage4_c49_s_fa3;
    wire stage4_c49_c_fa3;
    wire stage4_c50_s_fa0;
    wire stage4_c50_c_fa0;
    wire stage4_c50_s_fa1;
    wire stage4_c50_c_fa1;
    wire stage4_c50_s_fa2;
    wire stage4_c50_c_fa2;
    wire stage4_c50_s_fa3;
    wire stage4_c50_c_fa3;
    wire stage4_c51_s_fa0;
    wire stage4_c51_c_fa0;
    wire stage4_c51_s_fa1;
    wire stage4_c51_c_fa1;
    wire stage4_c51_s_fa2;
    wire stage4_c51_c_fa2;
    wire stage4_c51_s_fa3;
    wire stage4_c51_c_fa3;
    wire stage4_c52_s_fa0;
    wire stage4_c52_c_fa0;
    wire stage4_c52_s_fa1;
    wire stage4_c52_c_fa1;
    wire stage4_c52_s_fa2;
    wire stage4_c52_c_fa2;
    wire stage4_c52_s_fa3;
    wire stage4_c52_c_fa3;
    wire stage4_c53_s_fa0;
    wire stage4_c53_c_fa0;
    wire stage4_c53_s_fa1;
    wire stage4_c53_c_fa1;
    wire stage4_c53_s_fa2;
    wire stage4_c53_c_fa2;
    wire stage4_c53_s_fa3;
    wire stage4_c53_c_fa3;
    wire stage4_c54_s_fa0;
    wire stage4_c54_c_fa0;
    wire stage4_c54_s_fa1;
    wire stage4_c54_c_fa1;
    wire stage4_c54_s_fa2;
    wire stage4_c54_c_fa2;
    wire stage4_c54_s_fa3;
    wire stage4_c54_c_fa3;
    wire stage4_c55_s_fa0;
    wire stage4_c55_c_fa0;
    wire stage4_c55_s_fa1;
    wire stage4_c55_c_fa1;
    wire stage4_c55_s_fa2;
    wire stage4_c55_c_fa2;
    wire stage4_c55_s_fa3;
    wire stage4_c55_c_fa3;
    wire stage4_c56_s_fa0;
    wire stage4_c56_c_fa0;
    wire stage4_c56_s_fa1;
    wire stage4_c56_c_fa1;
    wire stage4_c56_s_fa2;
    wire stage4_c56_c_fa2;
    wire stage4_c56_s_fa3;
    wire stage4_c56_c_fa3;
    wire stage4_c57_s_fa0;
    wire stage4_c57_c_fa0;
    wire stage4_c57_s_fa1;
    wire stage4_c57_c_fa1;
    wire stage4_c57_s_fa2;
    wire stage4_c57_c_fa2;
    wire stage4_c57_s_fa3;
    wire stage4_c57_c_fa3;
    wire stage4_c58_s_fa0;
    wire stage4_c58_c_fa0;
    wire stage4_c58_s_fa1;
    wire stage4_c58_c_fa1;
    wire stage4_c58_s_fa2;
    wire stage4_c58_c_fa2;
    wire stage4_c58_s_fa3;
    wire stage4_c58_c_fa3;
    wire stage4_c59_s_fa0;
    wire stage4_c59_c_fa0;
    wire stage4_c59_s_fa1;
    wire stage4_c59_c_fa1;
    wire stage4_c59_s_fa2;
    wire stage4_c59_c_fa2;
    wire stage4_c59_s_fa3;
    wire stage4_c59_c_fa3;
    wire stage4_c60_s_fa0;
    wire stage4_c60_c_fa0;
    wire stage4_c60_s_fa1;
    wire stage4_c60_c_fa1;
    wire stage4_c60_s_fa2;
    wire stage4_c60_c_fa2;
    wire stage4_c60_s_fa3;
    wire stage4_c60_c_fa3;
    wire stage4_c61_s_fa0;
    wire stage4_c61_c_fa0;
    wire stage4_c61_s_fa1;
    wire stage4_c61_c_fa1;
    wire stage4_c61_s_fa2;
    wire stage4_c61_c_fa2;
    wire stage4_c61_s_fa3;
    wire stage4_c61_c_fa3;
    wire stage4_c62_s_fa0;
    wire stage4_c62_c_fa0;
    wire stage4_c62_s_fa1;
    wire stage4_c62_c_fa1;
    wire stage4_c62_s_fa2;
    wire stage4_c62_c_fa2;
    wire stage4_c62_s_fa3;
    wire stage4_c62_c_fa3;
    wire stage4_c63_s_fa0;
    wire stage4_c63_c_fa0;
    wire stage4_c63_s_fa1;
    wire stage4_c63_c_fa1;
    wire stage4_c63_s_fa2;
    wire stage4_c63_c_fa2;
    wire stage4_c63_s_fa3;
    wire stage4_c63_c_fa3;
    wire stage4_c64_s_fa0;
    wire stage4_c64_c_fa0;
    wire stage4_c64_s_fa1;
    wire stage4_c64_c_fa1;
    wire stage4_c64_s_fa2;
    wire stage4_c64_c_fa2;
    wire stage4_c64_s_fa3;
    wire stage4_c64_c_fa3;
    wire stage4_c65_s_fa0;
    wire stage4_c65_c_fa0;
    wire stage4_c65_s_fa1;
    wire stage4_c65_c_fa1;
    wire stage4_c65_s_fa2;
    wire stage4_c65_c_fa2;
    wire stage4_c65_s_fa3;
    wire stage4_c65_c_fa3;
    wire stage4_c66_s_fa0;
    wire stage4_c66_c_fa0;
    wire stage4_c66_s_fa1;
    wire stage4_c66_c_fa1;
    wire stage4_c66_s_fa2;
    wire stage4_c66_c_fa2;
    wire stage4_c66_s_fa3;
    wire stage4_c66_c_fa3;
    wire stage4_c67_s_fa0;
    wire stage4_c67_c_fa0;
    wire stage4_c67_s_fa1;
    wire stage4_c67_c_fa1;
    wire stage4_c67_s_fa2;
    wire stage4_c67_c_fa2;
    wire stage4_c67_s_fa3;
    wire stage4_c67_c_fa3;
    wire stage4_c68_s_fa0;
    wire stage4_c68_c_fa0;
    wire stage4_c68_s_fa1;
    wire stage4_c68_c_fa1;
    wire stage4_c68_s_fa2;
    wire stage4_c68_c_fa2;
    wire stage4_c68_s_fa3;
    wire stage4_c68_c_fa3;
    wire stage4_c69_s_fa0;
    wire stage4_c69_c_fa0;
    wire stage4_c69_s_fa1;
    wire stage4_c69_c_fa1;
    wire stage4_c69_s_fa2;
    wire stage4_c69_c_fa2;
    wire stage4_c69_s_fa3;
    wire stage4_c69_c_fa3;
    wire stage4_c70_s_fa0;
    wire stage4_c70_c_fa0;
    wire stage4_c70_s_fa1;
    wire stage4_c70_c_fa1;
    wire stage4_c70_s_fa2;
    wire stage4_c70_c_fa2;
    wire stage4_c70_s_fa3;
    wire stage4_c70_c_fa3;
    wire stage4_c71_s_fa0;
    wire stage4_c71_c_fa0;
    wire stage4_c71_s_fa1;
    wire stage4_c71_c_fa1;
    wire stage4_c71_s_fa2;
    wire stage4_c71_c_fa2;
    wire stage4_c71_s_fa3;
    wire stage4_c71_c_fa3;
    wire stage4_c72_s_fa0;
    wire stage4_c72_c_fa0;
    wire stage4_c72_s_fa1;
    wire stage4_c72_c_fa1;
    wire stage4_c72_s_fa2;
    wire stage4_c72_c_fa2;
    wire stage4_c72_s_fa3;
    wire stage4_c72_c_fa3;
    wire stage4_c73_s_fa0;
    wire stage4_c73_c_fa0;
    wire stage4_c73_s_fa1;
    wire stage4_c73_c_fa1;
    wire stage4_c73_s_fa2;
    wire stage4_c73_c_fa2;
    wire stage4_c73_s_fa3;
    wire stage4_c73_c_fa3;
    wire stage4_c74_s_fa0;
    wire stage4_c74_c_fa0;
    wire stage4_c74_s_fa1;
    wire stage4_c74_c_fa1;
    wire stage4_c74_s_fa2;
    wire stage4_c74_c_fa2;
    wire stage4_c74_s_fa3;
    wire stage4_c74_c_fa3;
    wire stage4_c75_s_fa0;
    wire stage4_c75_c_fa0;
    wire stage4_c75_s_fa1;
    wire stage4_c75_c_fa1;
    wire stage4_c75_s_fa2;
    wire stage4_c75_c_fa2;
    wire stage4_c75_s_fa3;
    wire stage4_c75_c_fa3;
    wire stage4_c76_s_fa0;
    wire stage4_c76_c_fa0;
    wire stage4_c76_s_fa1;
    wire stage4_c76_c_fa1;
    wire stage4_c76_s_fa2;
    wire stage4_c76_c_fa2;
    wire stage4_c76_s_fa3;
    wire stage4_c76_c_fa3;
    wire stage4_c77_s_fa0;
    wire stage4_c77_c_fa0;
    wire stage4_c77_s_fa1;
    wire stage4_c77_c_fa1;
    wire stage4_c77_s_fa2;
    wire stage4_c77_c_fa2;
    wire stage4_c77_s_fa3;
    wire stage4_c77_c_fa3;
    wire stage4_c78_s_fa0;
    wire stage4_c78_c_fa0;
    wire stage4_c78_s_fa1;
    wire stage4_c78_c_fa1;
    wire stage4_c78_s_fa2;
    wire stage4_c78_c_fa2;
    wire stage4_c78_s_ha0;
    wire stage4_c78_c_ha0;
    wire stage4_c79_s_fa0;
    wire stage4_c79_c_fa0;
    wire stage4_c79_s_fa1;
    wire stage4_c79_c_fa1;
    wire stage4_c79_s_fa2;
    wire stage4_c79_c_fa2;
    wire stage4_c79_s_ha0;
    wire stage4_c79_c_ha0;
    wire stage4_c80_s_fa0;
    wire stage4_c80_c_fa0;
    wire stage4_c80_s_fa1;
    wire stage4_c80_c_fa1;
    wire stage4_c80_s_fa2;
    wire stage4_c80_c_fa2;
    wire stage4_c81_s_fa0;
    wire stage4_c81_c_fa0;
    wire stage4_c81_s_fa1;
    wire stage4_c81_c_fa1;
    wire stage4_c81_s_fa2;
    wire stage4_c81_c_fa2;
    wire stage4_c82_s_fa0;
    wire stage4_c82_c_fa0;
    wire stage4_c82_s_fa1;
    wire stage4_c82_c_fa1;
    wire stage4_c82_s_fa2;
    wire stage4_c82_c_fa2;
    wire stage4_c83_s_fa0;
    wire stage4_c83_c_fa0;
    wire stage4_c83_s_fa1;
    wire stage4_c83_c_fa1;
    wire stage4_c83_s_fa2;
    wire stage4_c83_c_fa2;
    wire stage4_c84_s_fa0;
    wire stage4_c84_c_fa0;
    wire stage4_c84_s_fa1;
    wire stage4_c84_c_fa1;
    wire stage4_c84_s_fa2;
    wire stage4_c84_c_fa2;
    wire stage4_c85_s_fa0;
    wire stage4_c85_c_fa0;
    wire stage4_c85_s_fa1;
    wire stage4_c85_c_fa1;
    wire stage4_c85_s_fa2;
    wire stage4_c85_c_fa2;
    wire stage4_c86_s_fa0;
    wire stage4_c86_c_fa0;
    wire stage4_c86_s_fa1;
    wire stage4_c86_c_fa1;
    wire stage4_c86_s_ha0;
    wire stage4_c86_c_ha0;
    wire stage4_c87_s_fa0;
    wire stage4_c87_c_fa0;
    wire stage4_c87_s_fa1;
    wire stage4_c87_c_fa1;
    wire stage4_c87_s_ha0;
    wire stage4_c87_c_ha0;
    wire stage4_c88_s_fa0;
    wire stage4_c88_c_fa0;
    wire stage4_c88_s_fa1;
    wire stage4_c88_c_fa1;
    wire stage4_c88_s_ha0;
    wire stage4_c88_c_ha0;
    wire stage4_c89_s_fa0;
    wire stage4_c89_c_fa0;
    wire stage4_c89_s_fa1;
    wire stage4_c89_c_fa1;
    wire stage4_c89_s_ha0;
    wire stage4_c89_c_ha0;
    wire stage4_c90_s_fa0;
    wire stage4_c90_c_fa0;
    wire stage4_c90_s_fa1;
    wire stage4_c90_c_fa1;
    wire stage4_c90_s_ha0;
    wire stage4_c90_c_ha0;
    wire stage4_c91_s_fa0;
    wire stage4_c91_c_fa0;
    wire stage4_c91_s_fa1;
    wire stage4_c91_c_fa1;
    wire stage4_c91_s_ha0;
    wire stage4_c91_c_ha0;
    wire stage4_c92_s_fa0;
    wire stage4_c92_c_fa0;
    wire stage4_c92_s_fa1;
    wire stage4_c92_c_fa1;
    wire stage4_c93_s_fa0;
    wire stage4_c93_c_fa0;
    wire stage4_c93_s_fa1;
    wire stage4_c93_c_fa1;
    wire stage4_c94_s_fa0;
    wire stage4_c94_c_fa0;
    wire stage4_c94_s_fa1;
    wire stage4_c94_c_fa1;
    wire stage4_c95_s_fa0;
    wire stage4_c95_c_fa0;
    wire stage4_c95_s_fa1;
    wire stage4_c95_c_fa1;
    wire stage4_c96_s_fa0;
    wire stage4_c96_c_fa0;
    wire stage4_c96_s_fa1;
    wire stage4_c96_c_fa1;
    wire stage4_c97_s_fa0;
    wire stage4_c97_c_fa0;
    wire stage4_c97_s_fa1;
    wire stage4_c97_c_fa1;
    wire stage4_c98_s_fa0;
    wire stage4_c98_c_fa0;
    wire stage4_c98_s_fa1;
    wire stage4_c98_c_fa1;
    wire stage4_c99_s_fa0;
    wire stage4_c99_c_fa0;
    wire stage4_c99_s_ha0;
    wire stage4_c99_c_ha0;
    wire stage4_c100_s_fa0;
    wire stage4_c100_c_fa0;
    wire stage4_c101_s_fa0;
    wire stage4_c101_c_fa0;
    wire stage4_c102_s_fa0;
    wire stage4_c102_c_fa0;
    wire stage4_c103_s_fa0;
    wire stage4_c103_c_fa0;
    wire stage4_c104_s_fa0;
    wire stage4_c104_c_fa0;
    wire stage4_c105_s_fa0;
    wire stage4_c105_c_fa0;
    wire stage4_c106_s_fa0;
    wire stage4_c106_c_fa0;
    wire stage4_c107_s_ha0;
    wire stage4_c107_c_ha0;
    wire stage4_c108_s_ha0;
    wire stage4_c108_c_ha0;
    wire stage4_c109_s_ha0;
    wire stage4_c109_c_ha0;
    wire stage4_c110_s_ha0;
    wire stage4_c110_c_ha0;
    wire stage4_c111_s_ha0;
    wire stage4_c111_c_ha0;
    wire stage4_c112_s_ha0;
    wire stage4_c112_c_ha0;
    wire stage5_c5_s_ha0;
    wire stage5_c5_c_ha0;
    wire stage5_c6_s_ha0;
    wire stage5_c6_c_ha0;
    wire stage5_c7_s_ha0;
    wire stage5_c7_c_ha0;
    wire stage5_c8_s_ha0;
    wire stage5_c8_c_ha0;
    wire stage5_c9_s_ha0;
    wire stage5_c9_c_ha0;
    wire stage5_c10_s_fa0;
    wire stage5_c10_c_fa0;
    wire stage5_c11_s_fa0;
    wire stage5_c11_c_fa0;
    wire stage5_c12_s_fa0;
    wire stage5_c12_c_fa0;
    wire stage5_c13_s_fa0;
    wire stage5_c13_c_fa0;
    wire stage5_c14_s_fa0;
    wire stage5_c14_c_fa0;
    wire stage5_c15_s_fa0;
    wire stage5_c15_c_fa0;
    wire stage5_c16_s_fa0;
    wire stage5_c16_c_fa0;
    wire stage5_c17_s_fa0;
    wire stage5_c17_c_fa0;
    wire stage5_c18_s_fa0;
    wire stage5_c18_c_fa0;
    wire stage5_c19_s_fa0;
    wire stage5_c19_c_fa0;
    wire stage5_c20_s_fa0;
    wire stage5_c20_c_fa0;
    wire stage5_c21_s_fa0;
    wire stage5_c21_c_fa0;
    wire stage5_c21_s_ha0;
    wire stage5_c21_c_ha0;
    wire stage5_c22_s_fa0;
    wire stage5_c22_c_fa0;
    wire stage5_c22_s_ha0;
    wire stage5_c22_c_ha0;
    wire stage5_c23_s_fa0;
    wire stage5_c23_c_fa0;
    wire stage5_c23_s_ha0;
    wire stage5_c23_c_ha0;
    wire stage5_c24_s_fa0;
    wire stage5_c24_c_fa0;
    wire stage5_c24_s_ha0;
    wire stage5_c24_c_ha0;
    wire stage5_c25_s_fa0;
    wire stage5_c25_c_fa0;
    wire stage5_c25_s_fa1;
    wire stage5_c25_c_fa1;
    wire stage5_c26_s_fa0;
    wire stage5_c26_c_fa0;
    wire stage5_c26_s_fa1;
    wire stage5_c26_c_fa1;
    wire stage5_c27_s_fa0;
    wire stage5_c27_c_fa0;
    wire stage5_c27_s_fa1;
    wire stage5_c27_c_fa1;
    wire stage5_c28_s_fa0;
    wire stage5_c28_c_fa0;
    wire stage5_c28_s_fa1;
    wire stage5_c28_c_fa1;
    wire stage5_c29_s_fa0;
    wire stage5_c29_c_fa0;
    wire stage5_c29_s_fa1;
    wire stage5_c29_c_fa1;
    wire stage5_c30_s_fa0;
    wire stage5_c30_c_fa0;
    wire stage5_c30_s_fa1;
    wire stage5_c30_c_fa1;
    wire stage5_c31_s_fa0;
    wire stage5_c31_c_fa0;
    wire stage5_c31_s_fa1;
    wire stage5_c31_c_fa1;
    wire stage5_c32_s_fa0;
    wire stage5_c32_c_fa0;
    wire stage5_c32_s_fa1;
    wire stage5_c32_c_fa1;
    wire stage5_c33_s_fa0;
    wire stage5_c33_c_fa0;
    wire stage5_c33_s_fa1;
    wire stage5_c33_c_fa1;
    wire stage5_c34_s_fa0;
    wire stage5_c34_c_fa0;
    wire stage5_c34_s_fa1;
    wire stage5_c34_c_fa1;
    wire stage5_c35_s_fa0;
    wire stage5_c35_c_fa0;
    wire stage5_c35_s_fa1;
    wire stage5_c35_c_fa1;
    wire stage5_c35_s_ha0;
    wire stage5_c35_c_ha0;
    wire stage5_c36_s_fa0;
    wire stage5_c36_c_fa0;
    wire stage5_c36_s_fa1;
    wire stage5_c36_c_fa1;
    wire stage5_c36_s_ha0;
    wire stage5_c36_c_ha0;
    wire stage5_c37_s_fa0;
    wire stage5_c37_c_fa0;
    wire stage5_c37_s_fa1;
    wire stage5_c37_c_fa1;
    wire stage5_c37_s_ha0;
    wire stage5_c37_c_ha0;
    wire stage5_c38_s_fa0;
    wire stage5_c38_c_fa0;
    wire stage5_c38_s_fa1;
    wire stage5_c38_c_fa1;
    wire stage5_c38_s_ha0;
    wire stage5_c38_c_ha0;
    wire stage5_c39_s_fa0;
    wire stage5_c39_c_fa0;
    wire stage5_c39_s_fa1;
    wire stage5_c39_c_fa1;
    wire stage5_c39_s_ha0;
    wire stage5_c39_c_ha0;
    wire stage5_c40_s_fa0;
    wire stage5_c40_c_fa0;
    wire stage5_c40_s_fa1;
    wire stage5_c40_c_fa1;
    wire stage5_c40_s_ha0;
    wire stage5_c40_c_ha0;
    wire stage5_c41_s_fa0;
    wire stage5_c41_c_fa0;
    wire stage5_c41_s_fa1;
    wire stage5_c41_c_fa1;
    wire stage5_c41_s_fa2;
    wire stage5_c41_c_fa2;
    wire stage5_c42_s_fa0;
    wire stage5_c42_c_fa0;
    wire stage5_c42_s_fa1;
    wire stage5_c42_c_fa1;
    wire stage5_c42_s_fa2;
    wire stage5_c42_c_fa2;
    wire stage5_c43_s_fa0;
    wire stage5_c43_c_fa0;
    wire stage5_c43_s_fa1;
    wire stage5_c43_c_fa1;
    wire stage5_c43_s_fa2;
    wire stage5_c43_c_fa2;
    wire stage5_c44_s_fa0;
    wire stage5_c44_c_fa0;
    wire stage5_c44_s_fa1;
    wire stage5_c44_c_fa1;
    wire stage5_c44_s_fa2;
    wire stage5_c44_c_fa2;
    wire stage5_c45_s_fa0;
    wire stage5_c45_c_fa0;
    wire stage5_c45_s_fa1;
    wire stage5_c45_c_fa1;
    wire stage5_c45_s_fa2;
    wire stage5_c45_c_fa2;
    wire stage5_c46_s_fa0;
    wire stage5_c46_c_fa0;
    wire stage5_c46_s_fa1;
    wire stage5_c46_c_fa1;
    wire stage5_c46_s_fa2;
    wire stage5_c46_c_fa2;
    wire stage5_c47_s_fa0;
    wire stage5_c47_c_fa0;
    wire stage5_c47_s_fa1;
    wire stage5_c47_c_fa1;
    wire stage5_c47_s_fa2;
    wire stage5_c47_c_fa2;
    wire stage5_c48_s_fa0;
    wire stage5_c48_c_fa0;
    wire stage5_c48_s_fa1;
    wire stage5_c48_c_fa1;
    wire stage5_c48_s_fa2;
    wire stage5_c48_c_fa2;
    wire stage5_c49_s_fa0;
    wire stage5_c49_c_fa0;
    wire stage5_c49_s_fa1;
    wire stage5_c49_c_fa1;
    wire stage5_c49_s_fa2;
    wire stage5_c49_c_fa2;
    wire stage5_c50_s_fa0;
    wire stage5_c50_c_fa0;
    wire stage5_c50_s_fa1;
    wire stage5_c50_c_fa1;
    wire stage5_c50_s_fa2;
    wire stage5_c50_c_fa2;
    wire stage5_c51_s_fa0;
    wire stage5_c51_c_fa0;
    wire stage5_c51_s_fa1;
    wire stage5_c51_c_fa1;
    wire stage5_c51_s_fa2;
    wire stage5_c51_c_fa2;
    wire stage5_c52_s_fa0;
    wire stage5_c52_c_fa0;
    wire stage5_c52_s_fa1;
    wire stage5_c52_c_fa1;
    wire stage5_c52_s_fa2;
    wire stage5_c52_c_fa2;
    wire stage5_c53_s_fa0;
    wire stage5_c53_c_fa0;
    wire stage5_c53_s_fa1;
    wire stage5_c53_c_fa1;
    wire stage5_c53_s_fa2;
    wire stage5_c53_c_fa2;
    wire stage5_c54_s_fa0;
    wire stage5_c54_c_fa0;
    wire stage5_c54_s_fa1;
    wire stage5_c54_c_fa1;
    wire stage5_c54_s_fa2;
    wire stage5_c54_c_fa2;
    wire stage5_c55_s_fa0;
    wire stage5_c55_c_fa0;
    wire stage5_c55_s_fa1;
    wire stage5_c55_c_fa1;
    wire stage5_c55_s_fa2;
    wire stage5_c55_c_fa2;
    wire stage5_c56_s_fa0;
    wire stage5_c56_c_fa0;
    wire stage5_c56_s_fa1;
    wire stage5_c56_c_fa1;
    wire stage5_c56_s_fa2;
    wire stage5_c56_c_fa2;
    wire stage5_c57_s_fa0;
    wire stage5_c57_c_fa0;
    wire stage5_c57_s_fa1;
    wire stage5_c57_c_fa1;
    wire stage5_c57_s_fa2;
    wire stage5_c57_c_fa2;
    wire stage5_c58_s_fa0;
    wire stage5_c58_c_fa0;
    wire stage5_c58_s_fa1;
    wire stage5_c58_c_fa1;
    wire stage5_c58_s_fa2;
    wire stage5_c58_c_fa2;
    wire stage5_c59_s_fa0;
    wire stage5_c59_c_fa0;
    wire stage5_c59_s_fa1;
    wire stage5_c59_c_fa1;
    wire stage5_c59_s_fa2;
    wire stage5_c59_c_fa2;
    wire stage5_c60_s_fa0;
    wire stage5_c60_c_fa0;
    wire stage5_c60_s_fa1;
    wire stage5_c60_c_fa1;
    wire stage5_c60_s_fa2;
    wire stage5_c60_c_fa2;
    wire stage5_c61_s_fa0;
    wire stage5_c61_c_fa0;
    wire stage5_c61_s_fa1;
    wire stage5_c61_c_fa1;
    wire stage5_c61_s_fa2;
    wire stage5_c61_c_fa2;
    wire stage5_c62_s_fa0;
    wire stage5_c62_c_fa0;
    wire stage5_c62_s_fa1;
    wire stage5_c62_c_fa1;
    wire stage5_c62_s_fa2;
    wire stage5_c62_c_fa2;
    wire stage5_c63_s_fa0;
    wire stage5_c63_c_fa0;
    wire stage5_c63_s_fa1;
    wire stage5_c63_c_fa1;
    wire stage5_c63_s_fa2;
    wire stage5_c63_c_fa2;
    wire stage5_c64_s_fa0;
    wire stage5_c64_c_fa0;
    wire stage5_c64_s_fa1;
    wire stage5_c64_c_fa1;
    wire stage5_c64_s_fa2;
    wire stage5_c64_c_fa2;
    wire stage5_c65_s_fa0;
    wire stage5_c65_c_fa0;
    wire stage5_c65_s_fa1;
    wire stage5_c65_c_fa1;
    wire stage5_c65_s_fa2;
    wire stage5_c65_c_fa2;
    wire stage5_c66_s_fa0;
    wire stage5_c66_c_fa0;
    wire stage5_c66_s_fa1;
    wire stage5_c66_c_fa1;
    wire stage5_c66_s_fa2;
    wire stage5_c66_c_fa2;
    wire stage5_c67_s_fa0;
    wire stage5_c67_c_fa0;
    wire stage5_c67_s_fa1;
    wire stage5_c67_c_fa1;
    wire stage5_c67_s_fa2;
    wire stage5_c67_c_fa2;
    wire stage5_c68_s_fa0;
    wire stage5_c68_c_fa0;
    wire stage5_c68_s_fa1;
    wire stage5_c68_c_fa1;
    wire stage5_c68_s_fa2;
    wire stage5_c68_c_fa2;
    wire stage5_c69_s_fa0;
    wire stage5_c69_c_fa0;
    wire stage5_c69_s_fa1;
    wire stage5_c69_c_fa1;
    wire stage5_c69_s_fa2;
    wire stage5_c69_c_fa2;
    wire stage5_c70_s_fa0;
    wire stage5_c70_c_fa0;
    wire stage5_c70_s_fa1;
    wire stage5_c70_c_fa1;
    wire stage5_c70_s_fa2;
    wire stage5_c70_c_fa2;
    wire stage5_c71_s_fa0;
    wire stage5_c71_c_fa0;
    wire stage5_c71_s_fa1;
    wire stage5_c71_c_fa1;
    wire stage5_c71_s_fa2;
    wire stage5_c71_c_fa2;
    wire stage5_c72_s_fa0;
    wire stage5_c72_c_fa0;
    wire stage5_c72_s_fa1;
    wire stage5_c72_c_fa1;
    wire stage5_c72_s_fa2;
    wire stage5_c72_c_fa2;
    wire stage5_c73_s_fa0;
    wire stage5_c73_c_fa0;
    wire stage5_c73_s_fa1;
    wire stage5_c73_c_fa1;
    wire stage5_c73_s_ha0;
    wire stage5_c73_c_ha0;
    wire stage5_c74_s_fa0;
    wire stage5_c74_c_fa0;
    wire stage5_c74_s_fa1;
    wire stage5_c74_c_fa1;
    wire stage5_c74_s_ha0;
    wire stage5_c74_c_ha0;
    wire stage5_c75_s_fa0;
    wire stage5_c75_c_fa0;
    wire stage5_c75_s_fa1;
    wire stage5_c75_c_fa1;
    wire stage5_c75_s_ha0;
    wire stage5_c75_c_ha0;
    wire stage5_c76_s_fa0;
    wire stage5_c76_c_fa0;
    wire stage5_c76_s_fa1;
    wire stage5_c76_c_fa1;
    wire stage5_c76_s_ha0;
    wire stage5_c76_c_ha0;
    wire stage5_c77_s_fa0;
    wire stage5_c77_c_fa0;
    wire stage5_c77_s_fa1;
    wire stage5_c77_c_fa1;
    wire stage5_c77_s_ha0;
    wire stage5_c77_c_ha0;
    wire stage5_c78_s_fa0;
    wire stage5_c78_c_fa0;
    wire stage5_c78_s_fa1;
    wire stage5_c78_c_fa1;
    wire stage5_c78_s_ha0;
    wire stage5_c78_c_ha0;
    wire stage5_c79_s_fa0;
    wire stage5_c79_c_fa0;
    wire stage5_c79_s_fa1;
    wire stage5_c79_c_fa1;
    wire stage5_c79_s_ha0;
    wire stage5_c79_c_ha0;
    wire stage5_c80_s_fa0;
    wire stage5_c80_c_fa0;
    wire stage5_c80_s_fa1;
    wire stage5_c80_c_fa1;
    wire stage5_c80_s_ha0;
    wire stage5_c80_c_ha0;
    wire stage5_c81_s_fa0;
    wire stage5_c81_c_fa0;
    wire stage5_c81_s_fa1;
    wire stage5_c81_c_fa1;
    wire stage5_c82_s_fa0;
    wire stage5_c82_c_fa0;
    wire stage5_c82_s_fa1;
    wire stage5_c82_c_fa1;
    wire stage5_c83_s_fa0;
    wire stage5_c83_c_fa0;
    wire stage5_c83_s_fa1;
    wire stage5_c83_c_fa1;
    wire stage5_c84_s_fa0;
    wire stage5_c84_c_fa0;
    wire stage5_c84_s_fa1;
    wire stage5_c84_c_fa1;
    wire stage5_c85_s_fa0;
    wire stage5_c85_c_fa0;
    wire stage5_c85_s_fa1;
    wire stage5_c85_c_fa1;
    wire stage5_c86_s_fa0;
    wire stage5_c86_c_fa0;
    wire stage5_c86_s_fa1;
    wire stage5_c86_c_fa1;
    wire stage5_c87_s_fa0;
    wire stage5_c87_c_fa0;
    wire stage5_c87_s_fa1;
    wire stage5_c87_c_fa1;
    wire stage5_c88_s_fa0;
    wire stage5_c88_c_fa0;
    wire stage5_c88_s_fa1;
    wire stage5_c88_c_fa1;
    wire stage5_c89_s_fa0;
    wire stage5_c89_c_fa0;
    wire stage5_c89_s_fa1;
    wire stage5_c89_c_fa1;
    wire stage5_c90_s_fa0;
    wire stage5_c90_c_fa0;
    wire stage5_c90_s_fa1;
    wire stage5_c90_c_fa1;
    wire stage5_c91_s_fa0;
    wire stage5_c91_c_fa0;
    wire stage5_c91_s_fa1;
    wire stage5_c91_c_fa1;
    wire stage5_c92_s_fa0;
    wire stage5_c92_c_fa0;
    wire stage5_c92_s_fa1;
    wire stage5_c92_c_fa1;
    wire stage5_c93_s_fa0;
    wire stage5_c93_c_fa0;
    wire stage5_c93_s_ha0;
    wire stage5_c93_c_ha0;
    wire stage5_c94_s_fa0;
    wire stage5_c94_c_fa0;
    wire stage5_c95_s_fa0;
    wire stage5_c95_c_fa0;
    wire stage5_c96_s_fa0;
    wire stage5_c96_c_fa0;
    wire stage5_c97_s_fa0;
    wire stage5_c97_c_fa0;
    wire stage5_c98_s_fa0;
    wire stage5_c98_c_fa0;
    wire stage5_c99_s_fa0;
    wire stage5_c99_c_fa0;
    wire stage5_c100_s_fa0;
    wire stage5_c100_c_fa0;
    wire stage5_c101_s_fa0;
    wire stage5_c101_c_fa0;
    wire stage5_c102_s_fa0;
    wire stage5_c102_c_fa0;
    wire stage5_c103_s_fa0;
    wire stage5_c103_c_fa0;
    wire stage5_c104_s_fa0;
    wire stage5_c104_c_fa0;
    wire stage5_c105_s_ha0;
    wire stage5_c105_c_ha0;
    wire stage5_c106_s_ha0;
    wire stage5_c106_c_ha0;
    wire stage5_c107_s_ha0;
    wire stage5_c107_c_ha0;
    wire stage5_c108_s_ha0;
    wire stage5_c108_c_ha0;
    wire stage5_c109_s_ha0;
    wire stage5_c109_c_ha0;
    wire stage5_c110_s_ha0;
    wire stage5_c110_c_ha0;
    wire stage5_c111_s_ha0;
    wire stage5_c111_c_ha0;
    wire stage5_c112_s_ha0;
    wire stage5_c112_c_ha0;
    wire stage6_c6_s_ha0;
    wire stage6_c6_c_ha0;
    wire stage6_c7_s_ha0;
    wire stage6_c7_c_ha0;
    wire stage6_c8_s_ha0;
    wire stage6_c8_c_ha0;
    wire stage6_c9_s_ha0;
    wire stage6_c9_c_ha0;
    wire stage6_c10_s_ha0;
    wire stage6_c10_c_ha0;
    wire stage6_c11_s_ha0;
    wire stage6_c11_c_ha0;
    wire stage6_c12_s_ha0;
    wire stage6_c12_c_ha0;
    wire stage6_c13_s_ha0;
    wire stage6_c13_c_ha0;
    wire stage6_c14_s_ha0;
    wire stage6_c14_c_ha0;
    wire stage6_c15_s_fa0;
    wire stage6_c15_c_fa0;
    wire stage6_c16_s_fa0;
    wire stage6_c16_c_fa0;
    wire stage6_c17_s_fa0;
    wire stage6_c17_c_fa0;
    wire stage6_c18_s_fa0;
    wire stage6_c18_c_fa0;
    wire stage6_c19_s_fa0;
    wire stage6_c19_c_fa0;
    wire stage6_c20_s_fa0;
    wire stage6_c20_c_fa0;
    wire stage6_c21_s_fa0;
    wire stage6_c21_c_fa0;
    wire stage6_c22_s_fa0;
    wire stage6_c22_c_fa0;
    wire stage6_c23_s_fa0;
    wire stage6_c23_c_fa0;
    wire stage6_c24_s_fa0;
    wire stage6_c24_c_fa0;
    wire stage6_c25_s_fa0;
    wire stage6_c25_c_fa0;
    wire stage6_c26_s_fa0;
    wire stage6_c26_c_fa0;
    wire stage6_c27_s_fa0;
    wire stage6_c27_c_fa0;
    wire stage6_c28_s_fa0;
    wire stage6_c28_c_fa0;
    wire stage6_c29_s_fa0;
    wire stage6_c29_c_fa0;
    wire stage6_c30_s_fa0;
    wire stage6_c30_c_fa0;
    wire stage6_c31_s_fa0;
    wire stage6_c31_c_fa0;
    wire stage6_c31_s_ha0;
    wire stage6_c31_c_ha0;
    wire stage6_c32_s_fa0;
    wire stage6_c32_c_fa0;
    wire stage6_c32_s_ha0;
    wire stage6_c32_c_ha0;
    wire stage6_c33_s_fa0;
    wire stage6_c33_c_fa0;
    wire stage6_c33_s_ha0;
    wire stage6_c33_c_ha0;
    wire stage6_c34_s_fa0;
    wire stage6_c34_c_fa0;
    wire stage6_c34_s_ha0;
    wire stage6_c34_c_ha0;
    wire stage6_c35_s_fa0;
    wire stage6_c35_c_fa0;
    wire stage6_c35_s_ha0;
    wire stage6_c35_c_ha0;
    wire stage6_c36_s_fa0;
    wire stage6_c36_c_fa0;
    wire stage6_c36_s_fa1;
    wire stage6_c36_c_fa1;
    wire stage6_c37_s_fa0;
    wire stage6_c37_c_fa0;
    wire stage6_c37_s_fa1;
    wire stage6_c37_c_fa1;
    wire stage6_c38_s_fa0;
    wire stage6_c38_c_fa0;
    wire stage6_c38_s_fa1;
    wire stage6_c38_c_fa1;
    wire stage6_c39_s_fa0;
    wire stage6_c39_c_fa0;
    wire stage6_c39_s_fa1;
    wire stage6_c39_c_fa1;
    wire stage6_c40_s_fa0;
    wire stage6_c40_c_fa0;
    wire stage6_c40_s_fa1;
    wire stage6_c40_c_fa1;
    wire stage6_c41_s_fa0;
    wire stage6_c41_c_fa0;
    wire stage6_c41_s_fa1;
    wire stage6_c41_c_fa1;
    wire stage6_c42_s_fa0;
    wire stage6_c42_c_fa0;
    wire stage6_c42_s_fa1;
    wire stage6_c42_c_fa1;
    wire stage6_c43_s_fa0;
    wire stage6_c43_c_fa0;
    wire stage6_c43_s_fa1;
    wire stage6_c43_c_fa1;
    wire stage6_c44_s_fa0;
    wire stage6_c44_c_fa0;
    wire stage6_c44_s_fa1;
    wire stage6_c44_c_fa1;
    wire stage6_c45_s_fa0;
    wire stage6_c45_c_fa0;
    wire stage6_c45_s_fa1;
    wire stage6_c45_c_fa1;
    wire stage6_c46_s_fa0;
    wire stage6_c46_c_fa0;
    wire stage6_c46_s_fa1;
    wire stage6_c46_c_fa1;
    wire stage6_c47_s_fa0;
    wire stage6_c47_c_fa0;
    wire stage6_c47_s_fa1;
    wire stage6_c47_c_fa1;
    wire stage6_c48_s_fa0;
    wire stage6_c48_c_fa0;
    wire stage6_c48_s_fa1;
    wire stage6_c48_c_fa1;
    wire stage6_c49_s_fa0;
    wire stage6_c49_c_fa0;
    wire stage6_c49_s_fa1;
    wire stage6_c49_c_fa1;
    wire stage6_c50_s_fa0;
    wire stage6_c50_c_fa0;
    wire stage6_c50_s_fa1;
    wire stage6_c50_c_fa1;
    wire stage6_c51_s_fa0;
    wire stage6_c51_c_fa0;
    wire stage6_c51_s_fa1;
    wire stage6_c51_c_fa1;
    wire stage6_c52_s_fa0;
    wire stage6_c52_c_fa0;
    wire stage6_c52_s_fa1;
    wire stage6_c52_c_fa1;
    wire stage6_c53_s_fa0;
    wire stage6_c53_c_fa0;
    wire stage6_c53_s_fa1;
    wire stage6_c53_c_fa1;
    wire stage6_c54_s_fa0;
    wire stage6_c54_c_fa0;
    wire stage6_c54_s_fa1;
    wire stage6_c54_c_fa1;
    wire stage6_c55_s_fa0;
    wire stage6_c55_c_fa0;
    wire stage6_c55_s_fa1;
    wire stage6_c55_c_fa1;
    wire stage6_c56_s_fa0;
    wire stage6_c56_c_fa0;
    wire stage6_c56_s_fa1;
    wire stage6_c56_c_fa1;
    wire stage6_c57_s_fa0;
    wire stage6_c57_c_fa0;
    wire stage6_c57_s_fa1;
    wire stage6_c57_c_fa1;
    wire stage6_c58_s_fa0;
    wire stage6_c58_c_fa0;
    wire stage6_c58_s_fa1;
    wire stage6_c58_c_fa1;
    wire stage6_c59_s_fa0;
    wire stage6_c59_c_fa0;
    wire stage6_c59_s_fa1;
    wire stage6_c59_c_fa1;
    wire stage6_c60_s_fa0;
    wire stage6_c60_c_fa0;
    wire stage6_c60_s_fa1;
    wire stage6_c60_c_fa1;
    wire stage6_c61_s_fa0;
    wire stage6_c61_c_fa0;
    wire stage6_c61_s_fa1;
    wire stage6_c61_c_fa1;
    wire stage6_c62_s_fa0;
    wire stage6_c62_c_fa0;
    wire stage6_c62_s_fa1;
    wire stage6_c62_c_fa1;
    wire stage6_c63_s_fa0;
    wire stage6_c63_c_fa0;
    wire stage6_c63_s_fa1;
    wire stage6_c63_c_fa1;
    wire stage6_c64_s_fa0;
    wire stage6_c64_c_fa0;
    wire stage6_c64_s_fa1;
    wire stage6_c64_c_fa1;
    wire stage6_c65_s_fa0;
    wire stage6_c65_c_fa0;
    wire stage6_c65_s_fa1;
    wire stage6_c65_c_fa1;
    wire stage6_c66_s_fa0;
    wire stage6_c66_c_fa0;
    wire stage6_c66_s_fa1;
    wire stage6_c66_c_fa1;
    wire stage6_c67_s_fa0;
    wire stage6_c67_c_fa0;
    wire stage6_c67_s_fa1;
    wire stage6_c67_c_fa1;
    wire stage6_c68_s_fa0;
    wire stage6_c68_c_fa0;
    wire stage6_c68_s_fa1;
    wire stage6_c68_c_fa1;
    wire stage6_c69_s_fa0;
    wire stage6_c69_c_fa0;
    wire stage6_c69_s_fa1;
    wire stage6_c69_c_fa1;
    wire stage6_c70_s_fa0;
    wire stage6_c70_c_fa0;
    wire stage6_c70_s_fa1;
    wire stage6_c70_c_fa1;
    wire stage6_c71_s_fa0;
    wire stage6_c71_c_fa0;
    wire stage6_c71_s_fa1;
    wire stage6_c71_c_fa1;
    wire stage6_c72_s_fa0;
    wire stage6_c72_c_fa0;
    wire stage6_c72_s_fa1;
    wire stage6_c72_c_fa1;
    wire stage6_c73_s_fa0;
    wire stage6_c73_c_fa0;
    wire stage6_c73_s_fa1;
    wire stage6_c73_c_fa1;
    wire stage6_c74_s_fa0;
    wire stage6_c74_c_fa0;
    wire stage6_c74_s_fa1;
    wire stage6_c74_c_fa1;
    wire stage6_c75_s_fa0;
    wire stage6_c75_c_fa0;
    wire stage6_c75_s_fa1;
    wire stage6_c75_c_fa1;
    wire stage6_c76_s_fa0;
    wire stage6_c76_c_fa0;
    wire stage6_c76_s_fa1;
    wire stage6_c76_c_fa1;
    wire stage6_c77_s_fa0;
    wire stage6_c77_c_fa0;
    wire stage6_c77_s_fa1;
    wire stage6_c77_c_fa1;
    wire stage6_c78_s_fa0;
    wire stage6_c78_c_fa0;
    wire stage6_c78_s_fa1;
    wire stage6_c78_c_fa1;
    wire stage6_c79_s_fa0;
    wire stage6_c79_c_fa0;
    wire stage6_c79_s_fa1;
    wire stage6_c79_c_fa1;
    wire stage6_c80_s_fa0;
    wire stage6_c80_c_fa0;
    wire stage6_c80_s_fa1;
    wire stage6_c80_c_fa1;
    wire stage6_c81_s_fa0;
    wire stage6_c81_c_fa0;
    wire stage6_c81_s_fa1;
    wire stage6_c81_c_fa1;
    wire stage6_c82_s_fa0;
    wire stage6_c82_c_fa0;
    wire stage6_c82_s_ha0;
    wire stage6_c82_c_ha0;
    wire stage6_c83_s_fa0;
    wire stage6_c83_c_fa0;
    wire stage6_c83_s_ha0;
    wire stage6_c83_c_ha0;
    wire stage6_c84_s_fa0;
    wire stage6_c84_c_fa0;
    wire stage6_c84_s_ha0;
    wire stage6_c84_c_ha0;
    wire stage6_c85_s_fa0;
    wire stage6_c85_c_fa0;
    wire stage6_c85_s_ha0;
    wire stage6_c85_c_ha0;
    wire stage6_c86_s_fa0;
    wire stage6_c86_c_fa0;
    wire stage6_c87_s_fa0;
    wire stage6_c87_c_fa0;
    wire stage6_c88_s_fa0;
    wire stage6_c88_c_fa0;
    wire stage6_c89_s_fa0;
    wire stage6_c89_c_fa0;
    wire stage6_c90_s_fa0;
    wire stage6_c90_c_fa0;
    wire stage6_c91_s_fa0;
    wire stage6_c91_c_fa0;
    wire stage6_c92_s_fa0;
    wire stage6_c92_c_fa0;
    wire stage6_c93_s_fa0;
    wire stage6_c93_c_fa0;
    wire stage6_c94_s_fa0;
    wire stage6_c94_c_fa0;
    wire stage6_c95_s_fa0;
    wire stage6_c95_c_fa0;
    wire stage6_c96_s_fa0;
    wire stage6_c96_c_fa0;
    wire stage6_c97_s_fa0;
    wire stage6_c97_c_fa0;
    wire stage6_c98_s_fa0;
    wire stage6_c98_c_fa0;
    wire stage6_c99_s_fa0;
    wire stage6_c99_c_fa0;
    wire stage6_c100_s_fa0;
    wire stage6_c100_c_fa0;
    wire stage6_c101_s_ha0;
    wire stage6_c101_c_ha0;
    wire stage6_c102_s_ha0;
    wire stage6_c102_c_ha0;
    wire stage6_c103_s_ha0;
    wire stage6_c103_c_ha0;
    wire stage6_c104_s_ha0;
    wire stage6_c104_c_ha0;
    wire stage6_c105_s_ha0;
    wire stage6_c105_c_ha0;
    wire stage6_c106_s_ha0;
    wire stage6_c106_c_ha0;
    wire stage6_c107_s_ha0;
    wire stage6_c107_c_ha0;
    wire stage6_c108_s_ha0;
    wire stage6_c108_c_ha0;
    wire stage6_c109_s_ha0;
    wire stage6_c109_c_ha0;
    wire stage6_c110_s_ha0;
    wire stage6_c110_c_ha0;
    wire stage6_c111_s_ha0;
    wire stage6_c111_c_ha0;
    wire stage6_c112_s_ha0;
    wire stage6_c112_c_ha0;
    wire stage6_c113_s_ha0;
    wire stage6_c113_c_ha0;
    wire stage7_c7_s_ha0;
    wire stage7_c7_c_ha0;
    wire stage7_c8_s_ha0;
    wire stage7_c8_c_ha0;
    wire stage7_c9_s_ha0;
    wire stage7_c9_c_ha0;
    wire stage7_c10_s_ha0;
    wire stage7_c10_c_ha0;
    wire stage7_c11_s_ha0;
    wire stage7_c11_c_ha0;
    wire stage7_c12_s_ha0;
    wire stage7_c12_c_ha0;
    wire stage7_c13_s_ha0;
    wire stage7_c13_c_ha0;
    wire stage7_c14_s_ha0;
    wire stage7_c14_c_ha0;
    wire stage7_c15_s_ha0;
    wire stage7_c15_c_ha0;
    wire stage7_c16_s_ha0;
    wire stage7_c16_c_ha0;
    wire stage7_c17_s_ha0;
    wire stage7_c17_c_ha0;
    wire stage7_c18_s_ha0;
    wire stage7_c18_c_ha0;
    wire stage7_c19_s_ha0;
    wire stage7_c19_c_ha0;
    wire stage7_c20_s_ha0;
    wire stage7_c20_c_ha0;
    wire stage7_c21_s_ha0;
    wire stage7_c21_c_ha0;
    wire stage7_c22_s_fa0;
    wire stage7_c22_c_fa0;
    wire stage7_c23_s_fa0;
    wire stage7_c23_c_fa0;
    wire stage7_c24_s_fa0;
    wire stage7_c24_c_fa0;
    wire stage7_c25_s_fa0;
    wire stage7_c25_c_fa0;
    wire stage7_c26_s_fa0;
    wire stage7_c26_c_fa0;
    wire stage7_c27_s_fa0;
    wire stage7_c27_c_fa0;
    wire stage7_c28_s_fa0;
    wire stage7_c28_c_fa0;
    wire stage7_c29_s_fa0;
    wire stage7_c29_c_fa0;
    wire stage7_c30_s_fa0;
    wire stage7_c30_c_fa0;
    wire stage7_c31_s_fa0;
    wire stage7_c31_c_fa0;
    wire stage7_c32_s_fa0;
    wire stage7_c32_c_fa0;
    wire stage7_c33_s_fa0;
    wire stage7_c33_c_fa0;
    wire stage7_c34_s_fa0;
    wire stage7_c34_c_fa0;
    wire stage7_c35_s_fa0;
    wire stage7_c35_c_fa0;
    wire stage7_c36_s_fa0;
    wire stage7_c36_c_fa0;
    wire stage7_c37_s_fa0;
    wire stage7_c37_c_fa0;
    wire stage7_c38_s_fa0;
    wire stage7_c38_c_fa0;
    wire stage7_c39_s_fa0;
    wire stage7_c39_c_fa0;
    wire stage7_c40_s_fa0;
    wire stage7_c40_c_fa0;
    wire stage7_c41_s_fa0;
    wire stage7_c41_c_fa0;
    wire stage7_c42_s_fa0;
    wire stage7_c42_c_fa0;
    wire stage7_c43_s_fa0;
    wire stage7_c43_c_fa0;
    wire stage7_c44_s_fa0;
    wire stage7_c44_c_fa0;
    wire stage7_c45_s_fa0;
    wire stage7_c45_c_fa0;
    wire stage7_c46_s_fa0;
    wire stage7_c46_c_fa0;
    wire stage7_c47_s_fa0;
    wire stage7_c47_c_fa0;
    wire stage7_c48_s_fa0;
    wire stage7_c48_c_fa0;
    wire stage7_c49_s_fa0;
    wire stage7_c49_c_fa0;
    wire stage7_c50_s_fa0;
    wire stage7_c50_c_fa0;
    wire stage7_c51_s_fa0;
    wire stage7_c51_c_fa0;
    wire stage7_c52_s_fa0;
    wire stage7_c52_c_fa0;
    wire stage7_c53_s_fa0;
    wire stage7_c53_c_fa0;
    wire stage7_c54_s_fa0;
    wire stage7_c54_c_fa0;
    wire stage7_c55_s_fa0;
    wire stage7_c55_c_fa0;
    wire stage7_c56_s_fa0;
    wire stage7_c56_c_fa0;
    wire stage7_c57_s_fa0;
    wire stage7_c57_c_fa0;
    wire stage7_c58_s_fa0;
    wire stage7_c58_c_fa0;
    wire stage7_c59_s_fa0;
    wire stage7_c59_c_fa0;
    wire stage7_c60_s_fa0;
    wire stage7_c60_c_fa0;
    wire stage7_c61_s_fa0;
    wire stage7_c61_c_fa0;
    wire stage7_c62_s_fa0;
    wire stage7_c62_c_fa0;
    wire stage7_c63_s_fa0;
    wire stage7_c63_c_fa0;
    wire stage7_c64_s_fa0;
    wire stage7_c64_c_fa0;
    wire stage7_c65_s_fa0;
    wire stage7_c65_c_fa0;
    wire stage7_c66_s_fa0;
    wire stage7_c66_c_fa0;
    wire stage7_c67_s_fa0;
    wire stage7_c67_c_fa0;
    wire stage7_c68_s_fa0;
    wire stage7_c68_c_fa0;
    wire stage7_c69_s_fa0;
    wire stage7_c69_c_fa0;
    wire stage7_c70_s_fa0;
    wire stage7_c70_c_fa0;
    wire stage7_c71_s_fa0;
    wire stage7_c71_c_fa0;
    wire stage7_c72_s_fa0;
    wire stage7_c72_c_fa0;
    wire stage7_c73_s_fa0;
    wire stage7_c73_c_fa0;
    wire stage7_c74_s_fa0;
    wire stage7_c74_c_fa0;
    wire stage7_c75_s_fa0;
    wire stage7_c75_c_fa0;
    wire stage7_c76_s_fa0;
    wire stage7_c76_c_fa0;
    wire stage7_c77_s_fa0;
    wire stage7_c77_c_fa0;
    wire stage7_c78_s_fa0;
    wire stage7_c78_c_fa0;
    wire stage7_c79_s_fa0;
    wire stage7_c79_c_fa0;
    wire stage7_c80_s_fa0;
    wire stage7_c80_c_fa0;
    wire stage7_c81_s_fa0;
    wire stage7_c81_c_fa0;
    wire stage7_c82_s_fa0;
    wire stage7_c82_c_fa0;
    wire stage7_c83_s_fa0;
    wire stage7_c83_c_fa0;
    wire stage7_c84_s_fa0;
    wire stage7_c84_c_fa0;
    wire stage7_c85_s_fa0;
    wire stage7_c85_c_fa0;
    wire stage7_c86_s_fa0;
    wire stage7_c86_c_fa0;
    wire stage7_c87_s_fa0;
    wire stage7_c87_c_fa0;
    wire stage7_c88_s_fa0;
    wire stage7_c88_c_fa0;
    wire stage7_c89_s_fa0;
    wire stage7_c89_c_fa0;
    wire stage7_c90_s_fa0;
    wire stage7_c90_c_fa0;
    wire stage7_c91_s_fa0;
    wire stage7_c91_c_fa0;
    wire stage7_c92_s_fa0;
    wire stage7_c92_c_fa0;
    wire stage7_c93_s_fa0;
    wire stage7_c93_c_fa0;
    wire stage7_c94_s_fa0;
    wire stage7_c94_c_fa0;
    wire stage7_c95_s_ha0;
    wire stage7_c95_c_ha0;
    wire stage7_c96_s_ha0;
    wire stage7_c96_c_ha0;
    wire stage7_c97_s_ha0;
    wire stage7_c97_c_ha0;
    wire stage7_c98_s_ha0;
    wire stage7_c98_c_ha0;
    wire stage7_c99_s_ha0;
    wire stage7_c99_c_ha0;
    wire stage7_c100_s_ha0;
    wire stage7_c100_c_ha0;
    wire stage7_c101_s_ha0;
    wire stage7_c101_c_ha0;
    wire stage7_c102_s_ha0;
    wire stage7_c102_c_ha0;
    wire stage7_c103_s_ha0;
    wire stage7_c103_c_ha0;
    wire stage7_c104_s_ha0;
    wire stage7_c104_c_ha0;
    wire stage7_c105_s_ha0;
    wire stage7_c105_c_ha0;
    wire stage7_c106_s_ha0;
    wire stage7_c106_c_ha0;
    wire stage7_c107_s_ha0;
    wire stage7_c107_c_ha0;
    wire stage7_c108_s_ha0;
    wire stage7_c108_c_ha0;
    wire stage7_c109_s_ha0;
    wire stage7_c109_c_ha0;
    wire stage7_c110_s_ha0;
    wire stage7_c110_c_ha0;
    wire stage7_c111_s_ha0;
    wire stage7_c111_c_ha0;
    wire stage7_c112_s_ha0;
    wire stage7_c112_c_ha0;
    wire stage7_c113_s_ha0;
    wire stage7_c113_c_ha0;
    wire stage8_c8_s_ha0;
    wire stage8_c8_c_ha0;
    wire stage8_c9_s_ha0;
    wire stage8_c9_c_ha0;
    wire stage8_c10_s_ha0;
    wire stage8_c10_c_ha0;
    wire stage8_c11_s_ha0;
    wire stage8_c11_c_ha0;
    wire stage8_c12_s_ha0;
    wire stage8_c12_c_ha0;
    wire stage8_c13_s_ha0;
    wire stage8_c13_c_ha0;
    wire stage8_c14_s_ha0;
    wire stage8_c14_c_ha0;
    wire stage8_c15_s_ha0;
    wire stage8_c15_c_ha0;
    wire stage8_c16_s_ha0;
    wire stage8_c16_c_ha0;
    wire stage8_c17_s_ha0;
    wire stage8_c17_c_ha0;
    wire stage8_c18_s_ha0;
    wire stage8_c18_c_ha0;
    wire stage8_c19_s_ha0;
    wire stage8_c19_c_ha0;
    wire stage8_c20_s_ha0;
    wire stage8_c20_c_ha0;
    wire stage8_c21_s_ha0;
    wire stage8_c21_c_ha0;
    wire stage8_c22_s_ha0;
    wire stage8_c22_c_ha0;
    wire stage8_c23_s_ha0;
    wire stage8_c23_c_ha0;
    wire stage8_c24_s_ha0;
    wire stage8_c24_c_ha0;
    wire stage8_c25_s_ha0;
    wire stage8_c25_c_ha0;
    wire stage8_c26_s_ha0;
    wire stage8_c26_c_ha0;
    wire stage8_c27_s_ha0;
    wire stage8_c27_c_ha0;
    wire stage8_c28_s_ha0;
    wire stage8_c28_c_ha0;
    wire stage8_c29_s_ha0;
    wire stage8_c29_c_ha0;
    wire stage8_c30_s_ha0;
    wire stage8_c30_c_ha0;
    wire stage8_c31_s_ha0;
    wire stage8_c31_c_ha0;
    wire stage8_c32_s_fa0;
    wire stage8_c32_c_fa0;
    wire stage8_c33_s_fa0;
    wire stage8_c33_c_fa0;
    wire stage8_c34_s_fa0;
    wire stage8_c34_c_fa0;
    wire stage8_c35_s_fa0;
    wire stage8_c35_c_fa0;
    wire stage8_c36_s_fa0;
    wire stage8_c36_c_fa0;
    wire stage8_c37_s_fa0;
    wire stage8_c37_c_fa0;
    wire stage8_c38_s_fa0;
    wire stage8_c38_c_fa0;
    wire stage8_c39_s_fa0;
    wire stage8_c39_c_fa0;
    wire stage8_c40_s_fa0;
    wire stage8_c40_c_fa0;
    wire stage8_c41_s_fa0;
    wire stage8_c41_c_fa0;
    wire stage8_c42_s_fa0;
    wire stage8_c42_c_fa0;
    wire stage8_c43_s_fa0;
    wire stage8_c43_c_fa0;
    wire stage8_c44_s_fa0;
    wire stage8_c44_c_fa0;
    wire stage8_c45_s_fa0;
    wire stage8_c45_c_fa0;
    wire stage8_c46_s_fa0;
    wire stage8_c46_c_fa0;
    wire stage8_c47_s_fa0;
    wire stage8_c47_c_fa0;
    wire stage8_c48_s_fa0;
    wire stage8_c48_c_fa0;
    wire stage8_c49_s_fa0;
    wire stage8_c49_c_fa0;
    wire stage8_c50_s_fa0;
    wire stage8_c50_c_fa0;
    wire stage8_c51_s_fa0;
    wire stage8_c51_c_fa0;
    wire stage8_c52_s_fa0;
    wire stage8_c52_c_fa0;
    wire stage8_c53_s_fa0;
    wire stage8_c53_c_fa0;
    wire stage8_c54_s_fa0;
    wire stage8_c54_c_fa0;
    wire stage8_c55_s_fa0;
    wire stage8_c55_c_fa0;
    wire stage8_c56_s_fa0;
    wire stage8_c56_c_fa0;
    wire stage8_c57_s_fa0;
    wire stage8_c57_c_fa0;
    wire stage8_c58_s_fa0;
    wire stage8_c58_c_fa0;
    wire stage8_c59_s_fa0;
    wire stage8_c59_c_fa0;
    wire stage8_c60_s_fa0;
    wire stage8_c60_c_fa0;
    wire stage8_c61_s_fa0;
    wire stage8_c61_c_fa0;
    wire stage8_c62_s_fa0;
    wire stage8_c62_c_fa0;
    wire stage8_c63_s_fa0;
    wire stage8_c63_c_fa0;
    wire stage8_c64_s_fa0;
    wire stage8_c64_c_fa0;
    wire stage8_c65_s_fa0;
    wire stage8_c65_c_fa0;
    wire stage8_c66_s_fa0;
    wire stage8_c66_c_fa0;
    wire stage8_c67_s_fa0;
    wire stage8_c67_c_fa0;
    wire stage8_c68_s_fa0;
    wire stage8_c68_c_fa0;
    wire stage8_c69_s_fa0;
    wire stage8_c69_c_fa0;
    wire stage8_c70_s_fa0;
    wire stage8_c70_c_fa0;
    wire stage8_c71_s_fa0;
    wire stage8_c71_c_fa0;
    wire stage8_c72_s_fa0;
    wire stage8_c72_c_fa0;
    wire stage8_c73_s_fa0;
    wire stage8_c73_c_fa0;
    wire stage8_c74_s_fa0;
    wire stage8_c74_c_fa0;
    wire stage8_c75_s_fa0;
    wire stage8_c75_c_fa0;
    wire stage8_c76_s_fa0;
    wire stage8_c76_c_fa0;
    wire stage8_c77_s_fa0;
    wire stage8_c77_c_fa0;
    wire stage8_c78_s_fa0;
    wire stage8_c78_c_fa0;
    wire stage8_c79_s_fa0;
    wire stage8_c79_c_fa0;
    wire stage8_c80_s_fa0;
    wire stage8_c80_c_fa0;
    wire stage8_c81_s_fa0;
    wire stage8_c81_c_fa0;
    wire stage8_c82_s_fa0;
    wire stage8_c82_c_fa0;
    wire stage8_c83_s_fa0;
    wire stage8_c83_c_fa0;
    wire stage8_c84_s_fa0;
    wire stage8_c84_c_fa0;
    wire stage8_c85_s_fa0;
    wire stage8_c85_c_fa0;
    wire stage8_c86_s_fa0;
    wire stage8_c86_c_fa0;
    wire stage8_c87_s_ha0;
    wire stage8_c87_c_ha0;
    wire stage8_c88_s_ha0;
    wire stage8_c88_c_ha0;
    wire stage8_c89_s_ha0;
    wire stage8_c89_c_ha0;
    wire stage8_c90_s_ha0;
    wire stage8_c90_c_ha0;
    wire stage8_c91_s_ha0;
    wire stage8_c91_c_ha0;
    wire stage8_c92_s_ha0;
    wire stage8_c92_c_ha0;
    wire stage8_c93_s_ha0;
    wire stage8_c93_c_ha0;
    wire stage8_c94_s_ha0;
    wire stage8_c94_c_ha0;
    wire stage8_c95_s_ha0;
    wire stage8_c95_c_ha0;
    wire stage8_c96_s_ha0;
    wire stage8_c96_c_ha0;
    wire stage8_c97_s_ha0;
    wire stage8_c97_c_ha0;
    wire stage8_c98_s_ha0;
    wire stage8_c98_c_ha0;
    wire stage8_c99_s_ha0;
    wire stage8_c99_c_ha0;
    wire stage8_c100_s_ha0;
    wire stage8_c100_c_ha0;
    wire stage8_c101_s_ha0;
    wire stage8_c101_c_ha0;
    wire stage8_c102_s_ha0;
    wire stage8_c102_c_ha0;
    wire stage8_c103_s_ha0;
    wire stage8_c103_c_ha0;
    wire stage8_c104_s_ha0;
    wire stage8_c104_c_ha0;
    wire stage8_c105_s_ha0;
    wire stage8_c105_c_ha0;
    wire stage8_c106_s_ha0;
    wire stage8_c106_c_ha0;
    wire stage8_c107_s_ha0;
    wire stage8_c107_c_ha0;
    wire stage8_c108_s_ha0;
    wire stage8_c108_c_ha0;
    wire stage8_c109_s_ha0;
    wire stage8_c109_c_ha0;
    wire stage8_c110_s_ha0;
    wire stage8_c110_c_ha0;
    wire stage8_c111_s_ha0;
    wire stage8_c111_c_ha0;
    wire stage8_c112_s_ha0;
    wire stage8_c112_c_ha0;
    wire stage8_c113_s_ha0;
    wire stage8_c113_c_ha0;
    wire stage8_c114_s_ha0;
    wire stage8_c114_c_ha0;

    wire [112:0] final_add0 = {stage8_c114_c_ha0, stage8_c113_c_ha0, stage8_c112_c_ha0, stage8_c111_c_ha0, stage8_c110_c_ha0, stage8_c109_c_ha0, stage8_c108_c_ha0, stage8_c107_c_ha0, stage8_c106_c_ha0, stage8_c105_c_ha0, stage8_c104_c_ha0, stage8_c103_c_ha0, stage8_c102_c_ha0, stage8_c101_c_ha0, stage8_c100_c_ha0, stage8_c99_c_ha0, stage8_c98_c_ha0, stage8_c97_c_ha0, stage8_c96_c_ha0, stage8_c95_c_ha0, stage8_c94_c_ha0, stage8_c93_c_ha0, stage8_c92_c_ha0, stage8_c91_c_ha0, stage8_c90_c_ha0, stage8_c89_c_ha0, stage8_c88_c_ha0, stage8_c87_c_ha0, stage8_c86_c_fa0, stage8_c85_c_fa0, stage8_c84_c_fa0, stage8_c83_c_fa0, stage8_c82_c_fa0, stage8_c81_c_fa0, stage8_c80_c_fa0, stage8_c79_c_fa0, stage8_c78_c_fa0, stage8_c77_c_fa0, stage8_c76_c_fa0, stage8_c75_c_fa0, stage8_c74_c_fa0, stage8_c73_c_fa0, stage8_c72_c_fa0, stage8_c71_c_fa0, stage8_c70_c_fa0, stage8_c69_c_fa0, stage8_c68_c_fa0, stage8_c67_c_fa0, stage8_c66_c_fa0, stage8_c65_c_fa0, stage8_c64_c_fa0, stage8_c63_c_fa0, stage8_c62_c_fa0, stage8_c61_c_fa0, stage8_c60_c_fa0, stage8_c59_c_fa0, stage8_c58_c_fa0, stage8_c57_c_fa0, stage8_c56_c_fa0, stage8_c55_c_fa0, stage8_c54_c_fa0, stage8_c53_c_fa0, stage8_c52_c_fa0, stage8_c51_c_fa0, stage8_c50_c_fa0, stage8_c49_c_fa0, stage8_c48_c_fa0, stage8_c47_c_fa0, stage8_c46_c_fa0, stage8_c45_c_fa0, stage8_c44_c_fa0, stage8_c43_c_fa0, stage8_c42_c_fa0, stage8_c41_c_fa0, stage8_c40_c_fa0, stage8_c39_c_fa0, stage8_c38_c_fa0, stage8_c37_c_fa0, stage8_c36_c_fa0, stage8_c35_c_fa0, stage8_c34_c_fa0, stage8_c33_c_fa0, stage8_c32_c_fa0, stage8_c31_c_ha0, stage8_c30_c_ha0, stage8_c29_c_ha0, stage8_c28_c_ha0, stage8_c27_c_ha0, stage8_c26_c_ha0, stage8_c25_c_ha0, stage8_c24_c_ha0, stage8_c23_c_ha0, stage8_c22_c_ha0, stage8_c21_c_ha0, stage8_c20_c_ha0, stage8_c19_c_ha0, stage8_c18_c_ha0, stage8_c17_c_ha0, stage8_c16_c_ha0, stage8_c15_c_ha0, stage8_c14_c_ha0, stage8_c13_c_ha0, stage8_c12_c_ha0, stage8_c11_c_ha0, stage8_c10_c_ha0, stage8_c9_c_ha0, stage8_c8_c_ha0, stage8_c8_s_ha0, stage7_c7_s_ha0, stage6_c6_s_ha0, stage5_c5_s_ha0, stage4_c4_s_ha0, stage3_c3_s_ha0, stage2_c2_s_ha0, stage1_c1_s_ha0, stage0_r0_c0};

    wire [112:0] final_add1 = {1'b0, stage8_c114_s_ha0, stage8_c113_s_ha0, stage8_c112_s_ha0, stage8_c111_s_ha0, stage8_c110_s_ha0, stage8_c109_s_ha0, stage8_c108_s_ha0, stage8_c107_s_ha0, stage8_c106_s_ha0, stage8_c105_s_ha0, stage8_c104_s_ha0, stage8_c103_s_ha0, stage8_c102_s_ha0, stage8_c101_s_ha0, stage8_c100_s_ha0, stage8_c99_s_ha0, stage8_c98_s_ha0, stage8_c97_s_ha0, stage8_c96_s_ha0, stage8_c95_s_ha0, stage8_c94_s_ha0, stage8_c93_s_ha0, stage8_c92_s_ha0, stage8_c91_s_ha0, stage8_c90_s_ha0, stage8_c89_s_ha0, stage8_c88_s_ha0, stage8_c87_s_ha0, stage8_c86_s_fa0, stage8_c85_s_fa0, stage8_c84_s_fa0, stage8_c83_s_fa0, stage8_c82_s_fa0, stage8_c81_s_fa0, stage8_c80_s_fa0, stage8_c79_s_fa0, stage8_c78_s_fa0, stage8_c77_s_fa0, stage8_c76_s_fa0, stage8_c75_s_fa0, stage8_c74_s_fa0, stage8_c73_s_fa0, stage8_c72_s_fa0, stage8_c71_s_fa0, stage8_c70_s_fa0, stage8_c69_s_fa0, stage8_c68_s_fa0, stage8_c67_s_fa0, stage8_c66_s_fa0, stage8_c65_s_fa0, stage8_c64_s_fa0, stage8_c63_s_fa0, stage8_c62_s_fa0, stage8_c61_s_fa0, stage8_c60_s_fa0, stage8_c59_s_fa0, stage8_c58_s_fa0, stage8_c57_s_fa0, stage8_c56_s_fa0, stage8_c55_s_fa0, stage8_c54_s_fa0, stage8_c53_s_fa0, stage8_c52_s_fa0, stage8_c51_s_fa0, stage8_c50_s_fa0, stage8_c49_s_fa0, stage8_c48_s_fa0, stage8_c47_s_fa0, stage8_c46_s_fa0, stage8_c45_s_fa0, stage8_c44_s_fa0, stage8_c43_s_fa0, stage8_c42_s_fa0, stage8_c41_s_fa0, stage8_c40_s_fa0, stage8_c39_s_fa0, stage8_c38_s_fa0, stage8_c37_s_fa0, stage8_c36_s_fa0, stage8_c35_s_fa0, stage8_c34_s_fa0, stage8_c33_s_fa0, stage8_c32_s_fa0, stage8_c31_s_ha0, stage8_c30_s_ha0, stage8_c29_s_ha0, stage8_c28_s_ha0, stage8_c27_s_ha0, stage8_c26_s_ha0, stage8_c25_s_ha0, stage8_c24_s_ha0, stage8_c23_s_ha0, stage8_c22_s_ha0, stage8_c21_s_ha0, stage8_c20_s_ha0, stage8_c19_s_ha0, stage8_c18_s_ha0, stage8_c17_s_ha0, stage8_c16_s_ha0, stage8_c15_s_ha0, stage8_c14_s_ha0, stage8_c13_s_ha0, stage8_c12_s_ha0, stage8_c11_s_ha0, stage8_c10_s_ha0, stage8_c9_s_ha0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};

    assign P = final_add0 + final_add1;
    //the logic
    assign stage0_r0_c0 = A[0] & B[0];
    assign stage0_r0_c1 = A[0] & B[1];
    assign stage0_r1_c0 = A[1] & B[0];
    assign stage0_r0_c2 = A[0] & B[2];
    assign stage0_r1_c1 = A[1] & B[1];
    assign stage0_r2_c0 = A[2] & B[0];
    assign stage0_r0_c3 = A[0] & B[3];
    assign stage0_r1_c2 = A[1] & B[2];
    assign stage0_r2_c1 = A[2] & B[1];
    assign stage0_r3_c0 = A[3] & B[0];
    assign stage0_r0_c4 = A[0] & B[4];
    assign stage0_r1_c3 = A[1] & B[3];
    assign stage0_r2_c2 = A[2] & B[2];
    assign stage0_r3_c1 = A[3] & B[1];
    assign stage0_r4_c0 = A[4] & B[0];
    assign stage0_r0_c5 = A[0] & B[5];
    assign stage0_r1_c4 = A[1] & B[4];
    assign stage0_r2_c3 = A[2] & B[3];
    assign stage0_r3_c2 = A[3] & B[2];
    assign stage0_r4_c1 = A[4] & B[1];
    assign stage0_r5_c0 = A[5] & B[0];
    assign stage0_r0_c6 = A[0] & B[6];
    assign stage0_r1_c5 = A[1] & B[5];
    assign stage0_r2_c4 = A[2] & B[4];
    assign stage0_r3_c3 = A[3] & B[3];
    assign stage0_r4_c2 = A[4] & B[2];
    assign stage0_r5_c1 = A[5] & B[1];
    assign stage0_r6_c0 = A[6] & B[0];
    assign stage0_r0_c7 = A[0] & B[7];
    assign stage0_r1_c6 = A[1] & B[6];
    assign stage0_r2_c5 = A[2] & B[5];
    assign stage0_r3_c4 = A[3] & B[4];
    assign stage0_r4_c3 = A[4] & B[3];
    assign stage0_r5_c2 = A[5] & B[2];
    assign stage0_r6_c1 = A[6] & B[1];
    assign stage0_r7_c0 = A[7] & B[0];
    assign stage0_r0_c8 = A[0] & B[8];
    assign stage0_r1_c7 = A[1] & B[7];
    assign stage0_r2_c6 = A[2] & B[6];
    assign stage0_r3_c5 = A[3] & B[5];
    assign stage0_r4_c4 = A[4] & B[4];
    assign stage0_r5_c3 = A[5] & B[3];
    assign stage0_r6_c2 = A[6] & B[2];
    assign stage0_r7_c1 = A[7] & B[1];
    assign stage0_r8_c0 = A[8] & B[0];
    assign stage0_r0_c9 = A[0] & B[9];
    assign stage0_r1_c8 = A[1] & B[8];
    assign stage0_r2_c7 = A[2] & B[7];
    assign stage0_r3_c6 = A[3] & B[6];
    assign stage0_r4_c5 = A[4] & B[5];
    assign stage0_r5_c4 = A[5] & B[4];
    assign stage0_r6_c3 = A[6] & B[3];
    assign stage0_r7_c2 = A[7] & B[2];
    assign stage0_r8_c1 = A[8] & B[1];
    assign stage0_r9_c0 = A[9] & B[0];
    assign stage0_r0_c10 = A[0] & B[10];
    assign stage0_r1_c9 = A[1] & B[9];
    assign stage0_r2_c8 = A[2] & B[8];
    assign stage0_r3_c7 = A[3] & B[7];
    assign stage0_r4_c6 = A[4] & B[6];
    assign stage0_r5_c5 = A[5] & B[5];
    assign stage0_r6_c4 = A[6] & B[4];
    assign stage0_r7_c3 = A[7] & B[3];
    assign stage0_r8_c2 = A[8] & B[2];
    assign stage0_r9_c1 = A[9] & B[1];
    assign stage0_r10_c0 = A[10] & B[0];
    assign stage0_r0_c11 = A[0] & B[11];
    assign stage0_r1_c10 = A[1] & B[10];
    assign stage0_r2_c9 = A[2] & B[9];
    assign stage0_r3_c8 = A[3] & B[8];
    assign stage0_r4_c7 = A[4] & B[7];
    assign stage0_r5_c6 = A[5] & B[6];
    assign stage0_r6_c5 = A[6] & B[5];
    assign stage0_r7_c4 = A[7] & B[4];
    assign stage0_r8_c3 = A[8] & B[3];
    assign stage0_r9_c2 = A[9] & B[2];
    assign stage0_r10_c1 = A[10] & B[1];
    assign stage0_r11_c0 = A[11] & B[0];
    assign stage0_r0_c12 = A[0] & B[12];
    assign stage0_r1_c11 = A[1] & B[11];
    assign stage0_r2_c10 = A[2] & B[10];
    assign stage0_r3_c9 = A[3] & B[9];
    assign stage0_r4_c8 = A[4] & B[8];
    assign stage0_r5_c7 = A[5] & B[7];
    assign stage0_r6_c6 = A[6] & B[6];
    assign stage0_r7_c5 = A[7] & B[5];
    assign stage0_r8_c4 = A[8] & B[4];
    assign stage0_r9_c3 = A[9] & B[3];
    assign stage0_r10_c2 = A[10] & B[2];
    assign stage0_r11_c1 = A[11] & B[1];
    assign stage0_r12_c0 = A[12] & B[0];
    assign stage0_r0_c13 = A[0] & B[13];
    assign stage0_r1_c12 = A[1] & B[12];
    assign stage0_r2_c11 = A[2] & B[11];
    assign stage0_r3_c10 = A[3] & B[10];
    assign stage0_r4_c9 = A[4] & B[9];
    assign stage0_r5_c8 = A[5] & B[8];
    assign stage0_r6_c7 = A[6] & B[7];
    assign stage0_r7_c6 = A[7] & B[6];
    assign stage0_r8_c5 = A[8] & B[5];
    assign stage0_r9_c4 = A[9] & B[4];
    assign stage0_r10_c3 = A[10] & B[3];
    assign stage0_r11_c2 = A[11] & B[2];
    assign stage0_r12_c1 = A[12] & B[1];
    assign stage0_r13_c0 = A[13] & B[0];
    assign stage0_r0_c14 = A[0] & B[14];
    assign stage0_r1_c13 = A[1] & B[13];
    assign stage0_r2_c12 = A[2] & B[12];
    assign stage0_r3_c11 = A[3] & B[11];
    assign stage0_r4_c10 = A[4] & B[10];
    assign stage0_r5_c9 = A[5] & B[9];
    assign stage0_r6_c8 = A[6] & B[8];
    assign stage0_r7_c7 = A[7] & B[7];
    assign stage0_r8_c6 = A[8] & B[6];
    assign stage0_r9_c5 = A[9] & B[5];
    assign stage0_r10_c4 = A[10] & B[4];
    assign stage0_r11_c3 = A[11] & B[3];
    assign stage0_r12_c2 = A[12] & B[2];
    assign stage0_r13_c1 = A[13] & B[1];
    assign stage0_r14_c0 = A[14] & B[0];
    assign stage0_r0_c15 = A[0] & B[15];
    assign stage0_r1_c14 = A[1] & B[14];
    assign stage0_r2_c13 = A[2] & B[13];
    assign stage0_r3_c12 = A[3] & B[12];
    assign stage0_r4_c11 = A[4] & B[11];
    assign stage0_r5_c10 = A[5] & B[10];
    assign stage0_r6_c9 = A[6] & B[9];
    assign stage0_r7_c8 = A[7] & B[8];
    assign stage0_r8_c7 = A[8] & B[7];
    assign stage0_r9_c6 = A[9] & B[6];
    assign stage0_r10_c5 = A[10] & B[5];
    assign stage0_r11_c4 = A[11] & B[4];
    assign stage0_r12_c3 = A[12] & B[3];
    assign stage0_r13_c2 = A[13] & B[2];
    assign stage0_r14_c1 = A[14] & B[1];
    assign stage0_r15_c0 = A[15] & B[0];
    assign stage0_r0_c16 = A[0] & B[16];
    assign stage0_r1_c15 = A[1] & B[15];
    assign stage0_r2_c14 = A[2] & B[14];
    assign stage0_r3_c13 = A[3] & B[13];
    assign stage0_r4_c12 = A[4] & B[12];
    assign stage0_r5_c11 = A[5] & B[11];
    assign stage0_r6_c10 = A[6] & B[10];
    assign stage0_r7_c9 = A[7] & B[9];
    assign stage0_r8_c8 = A[8] & B[8];
    assign stage0_r9_c7 = A[9] & B[7];
    assign stage0_r10_c6 = A[10] & B[6];
    assign stage0_r11_c5 = A[11] & B[5];
    assign stage0_r12_c4 = A[12] & B[4];
    assign stage0_r13_c3 = A[13] & B[3];
    assign stage0_r14_c2 = A[14] & B[2];
    assign stage0_r15_c1 = A[15] & B[1];
    assign stage0_r16_c0 = A[16] & B[0];
    assign stage0_r0_c17 = A[0] & B[17];
    assign stage0_r1_c16 = A[1] & B[16];
    assign stage0_r2_c15 = A[2] & B[15];
    assign stage0_r3_c14 = A[3] & B[14];
    assign stage0_r4_c13 = A[4] & B[13];
    assign stage0_r5_c12 = A[5] & B[12];
    assign stage0_r6_c11 = A[6] & B[11];
    assign stage0_r7_c10 = A[7] & B[10];
    assign stage0_r8_c9 = A[8] & B[9];
    assign stage0_r9_c8 = A[9] & B[8];
    assign stage0_r10_c7 = A[10] & B[7];
    assign stage0_r11_c6 = A[11] & B[6];
    assign stage0_r12_c5 = A[12] & B[5];
    assign stage0_r13_c4 = A[13] & B[4];
    assign stage0_r14_c3 = A[14] & B[3];
    assign stage0_r15_c2 = A[15] & B[2];
    assign stage0_r16_c1 = A[16] & B[1];
    assign stage0_r17_c0 = A[17] & B[0];
    assign stage0_r0_c18 = A[0] & B[18];
    assign stage0_r1_c17 = A[1] & B[17];
    assign stage0_r2_c16 = A[2] & B[16];
    assign stage0_r3_c15 = A[3] & B[15];
    assign stage0_r4_c14 = A[4] & B[14];
    assign stage0_r5_c13 = A[5] & B[13];
    assign stage0_r6_c12 = A[6] & B[12];
    assign stage0_r7_c11 = A[7] & B[11];
    assign stage0_r8_c10 = A[8] & B[10];
    assign stage0_r9_c9 = A[9] & B[9];
    assign stage0_r10_c8 = A[10] & B[8];
    assign stage0_r11_c7 = A[11] & B[7];
    assign stage0_r12_c6 = A[12] & B[6];
    assign stage0_r13_c5 = A[13] & B[5];
    assign stage0_r14_c4 = A[14] & B[4];
    assign stage0_r15_c3 = A[15] & B[3];
    assign stage0_r16_c2 = A[16] & B[2];
    assign stage0_r17_c1 = A[17] & B[1];
    assign stage0_r18_c0 = A[18] & B[0];
    assign stage0_r0_c19 = A[0] & B[19];
    assign stage0_r1_c18 = A[1] & B[18];
    assign stage0_r2_c17 = A[2] & B[17];
    assign stage0_r3_c16 = A[3] & B[16];
    assign stage0_r4_c15 = A[4] & B[15];
    assign stage0_r5_c14 = A[5] & B[14];
    assign stage0_r6_c13 = A[6] & B[13];
    assign stage0_r7_c12 = A[7] & B[12];
    assign stage0_r8_c11 = A[8] & B[11];
    assign stage0_r9_c10 = A[9] & B[10];
    assign stage0_r10_c9 = A[10] & B[9];
    assign stage0_r11_c8 = A[11] & B[8];
    assign stage0_r12_c7 = A[12] & B[7];
    assign stage0_r13_c6 = A[13] & B[6];
    assign stage0_r14_c5 = A[14] & B[5];
    assign stage0_r15_c4 = A[15] & B[4];
    assign stage0_r16_c3 = A[16] & B[3];
    assign stage0_r17_c2 = A[17] & B[2];
    assign stage0_r18_c1 = A[18] & B[1];
    assign stage0_r19_c0 = A[19] & B[0];
    assign stage0_r0_c20 = A[0] & B[20];
    assign stage0_r1_c19 = A[1] & B[19];
    assign stage0_r2_c18 = A[2] & B[18];
    assign stage0_r3_c17 = A[3] & B[17];
    assign stage0_r4_c16 = A[4] & B[16];
    assign stage0_r5_c15 = A[5] & B[15];
    assign stage0_r6_c14 = A[6] & B[14];
    assign stage0_r7_c13 = A[7] & B[13];
    assign stage0_r8_c12 = A[8] & B[12];
    assign stage0_r9_c11 = A[9] & B[11];
    assign stage0_r10_c10 = A[10] & B[10];
    assign stage0_r11_c9 = A[11] & B[9];
    assign stage0_r12_c8 = A[12] & B[8];
    assign stage0_r13_c7 = A[13] & B[7];
    assign stage0_r14_c6 = A[14] & B[6];
    assign stage0_r15_c5 = A[15] & B[5];
    assign stage0_r16_c4 = A[16] & B[4];
    assign stage0_r17_c3 = A[17] & B[3];
    assign stage0_r18_c2 = A[18] & B[2];
    assign stage0_r19_c1 = A[19] & B[1];
    assign stage0_r20_c0 = A[20] & B[0];
    assign stage0_r0_c21 = A[0] & B[21];
    assign stage0_r1_c20 = A[1] & B[20];
    assign stage0_r2_c19 = A[2] & B[19];
    assign stage0_r3_c18 = A[3] & B[18];
    assign stage0_r4_c17 = A[4] & B[17];
    assign stage0_r5_c16 = A[5] & B[16];
    assign stage0_r6_c15 = A[6] & B[15];
    assign stage0_r7_c14 = A[7] & B[14];
    assign stage0_r8_c13 = A[8] & B[13];
    assign stage0_r9_c12 = A[9] & B[12];
    assign stage0_r10_c11 = A[10] & B[11];
    assign stage0_r11_c10 = A[11] & B[10];
    assign stage0_r12_c9 = A[12] & B[9];
    assign stage0_r13_c8 = A[13] & B[8];
    assign stage0_r14_c7 = A[14] & B[7];
    assign stage0_r15_c6 = A[15] & B[6];
    assign stage0_r16_c5 = A[16] & B[5];
    assign stage0_r17_c4 = A[17] & B[4];
    assign stage0_r18_c3 = A[18] & B[3];
    assign stage0_r19_c2 = A[19] & B[2];
    assign stage0_r20_c1 = A[20] & B[1];
    assign stage0_r21_c0 = A[21] & B[0];
    assign stage0_r0_c22 = A[0] & B[22];
    assign stage0_r1_c21 = A[1] & B[21];
    assign stage0_r2_c20 = A[2] & B[20];
    assign stage0_r3_c19 = A[3] & B[19];
    assign stage0_r4_c18 = A[4] & B[18];
    assign stage0_r5_c17 = A[5] & B[17];
    assign stage0_r6_c16 = A[6] & B[16];
    assign stage0_r7_c15 = A[7] & B[15];
    assign stage0_r8_c14 = A[8] & B[14];
    assign stage0_r9_c13 = A[9] & B[13];
    assign stage0_r10_c12 = A[10] & B[12];
    assign stage0_r11_c11 = A[11] & B[11];
    assign stage0_r12_c10 = A[12] & B[10];
    assign stage0_r13_c9 = A[13] & B[9];
    assign stage0_r14_c8 = A[14] & B[8];
    assign stage0_r15_c7 = A[15] & B[7];
    assign stage0_r16_c6 = A[16] & B[6];
    assign stage0_r17_c5 = A[17] & B[5];
    assign stage0_r18_c4 = A[18] & B[4];
    assign stage0_r19_c3 = A[19] & B[3];
    assign stage0_r20_c2 = A[20] & B[2];
    assign stage0_r21_c1 = A[21] & B[1];
    assign stage0_r22_c0 = A[22] & B[0];
    assign stage0_r0_c23 = A[0] & B[23];
    assign stage0_r1_c22 = A[1] & B[22];
    assign stage0_r2_c21 = A[2] & B[21];
    assign stage0_r3_c20 = A[3] & B[20];
    assign stage0_r4_c19 = A[4] & B[19];
    assign stage0_r5_c18 = A[5] & B[18];
    assign stage0_r6_c17 = A[6] & B[17];
    assign stage0_r7_c16 = A[7] & B[16];
    assign stage0_r8_c15 = A[8] & B[15];
    assign stage0_r9_c14 = A[9] & B[14];
    assign stage0_r10_c13 = A[10] & B[13];
    assign stage0_r11_c12 = A[11] & B[12];
    assign stage0_r12_c11 = A[12] & B[11];
    assign stage0_r13_c10 = A[13] & B[10];
    assign stage0_r14_c9 = A[14] & B[9];
    assign stage0_r15_c8 = A[15] & B[8];
    assign stage0_r16_c7 = A[16] & B[7];
    assign stage0_r17_c6 = A[17] & B[6];
    assign stage0_r18_c5 = A[18] & B[5];
    assign stage0_r19_c4 = A[19] & B[4];
    assign stage0_r20_c3 = A[20] & B[3];
    assign stage0_r21_c2 = A[21] & B[2];
    assign stage0_r22_c1 = A[22] & B[1];
    assign stage0_r23_c0 = A[23] & B[0];
    assign stage0_r0_c24 = A[0] & B[24];
    assign stage0_r1_c23 = A[1] & B[23];
    assign stage0_r2_c22 = A[2] & B[22];
    assign stage0_r3_c21 = A[3] & B[21];
    assign stage0_r4_c20 = A[4] & B[20];
    assign stage0_r5_c19 = A[5] & B[19];
    assign stage0_r6_c18 = A[6] & B[18];
    assign stage0_r7_c17 = A[7] & B[17];
    assign stage0_r8_c16 = A[8] & B[16];
    assign stage0_r9_c15 = A[9] & B[15];
    assign stage0_r10_c14 = A[10] & B[14];
    assign stage0_r11_c13 = A[11] & B[13];
    assign stage0_r12_c12 = A[12] & B[12];
    assign stage0_r13_c11 = A[13] & B[11];
    assign stage0_r14_c10 = A[14] & B[10];
    assign stage0_r15_c9 = A[15] & B[9];
    assign stage0_r16_c8 = A[16] & B[8];
    assign stage0_r17_c7 = A[17] & B[7];
    assign stage0_r18_c6 = A[18] & B[6];
    assign stage0_r19_c5 = A[19] & B[5];
    assign stage0_r20_c4 = A[20] & B[4];
    assign stage0_r21_c3 = A[21] & B[3];
    assign stage0_r22_c2 = A[22] & B[2];
    assign stage0_r23_c1 = A[23] & B[1];
    assign stage0_r24_c0 = A[24] & B[0];
    assign stage0_r0_c25 = A[0] & B[25];
    assign stage0_r1_c24 = A[1] & B[24];
    assign stage0_r2_c23 = A[2] & B[23];
    assign stage0_r3_c22 = A[3] & B[22];
    assign stage0_r4_c21 = A[4] & B[21];
    assign stage0_r5_c20 = A[5] & B[20];
    assign stage0_r6_c19 = A[6] & B[19];
    assign stage0_r7_c18 = A[7] & B[18];
    assign stage0_r8_c17 = A[8] & B[17];
    assign stage0_r9_c16 = A[9] & B[16];
    assign stage0_r10_c15 = A[10] & B[15];
    assign stage0_r11_c14 = A[11] & B[14];
    assign stage0_r12_c13 = A[12] & B[13];
    assign stage0_r13_c12 = A[13] & B[12];
    assign stage0_r14_c11 = A[14] & B[11];
    assign stage0_r15_c10 = A[15] & B[10];
    assign stage0_r16_c9 = A[16] & B[9];
    assign stage0_r17_c8 = A[17] & B[8];
    assign stage0_r18_c7 = A[18] & B[7];
    assign stage0_r19_c6 = A[19] & B[6];
    assign stage0_r20_c5 = A[20] & B[5];
    assign stage0_r21_c4 = A[21] & B[4];
    assign stage0_r22_c3 = A[22] & B[3];
    assign stage0_r23_c2 = A[23] & B[2];
    assign stage0_r24_c1 = A[24] & B[1];
    assign stage0_r25_c0 = A[25] & B[0];
    assign stage0_r0_c26 = A[0] & B[26];
    assign stage0_r1_c25 = A[1] & B[25];
    assign stage0_r2_c24 = A[2] & B[24];
    assign stage0_r3_c23 = A[3] & B[23];
    assign stage0_r4_c22 = A[4] & B[22];
    assign stage0_r5_c21 = A[5] & B[21];
    assign stage0_r6_c20 = A[6] & B[20];
    assign stage0_r7_c19 = A[7] & B[19];
    assign stage0_r8_c18 = A[8] & B[18];
    assign stage0_r9_c17 = A[9] & B[17];
    assign stage0_r10_c16 = A[10] & B[16];
    assign stage0_r11_c15 = A[11] & B[15];
    assign stage0_r12_c14 = A[12] & B[14];
    assign stage0_r13_c13 = A[13] & B[13];
    assign stage0_r14_c12 = A[14] & B[12];
    assign stage0_r15_c11 = A[15] & B[11];
    assign stage0_r16_c10 = A[16] & B[10];
    assign stage0_r17_c9 = A[17] & B[9];
    assign stage0_r18_c8 = A[18] & B[8];
    assign stage0_r19_c7 = A[19] & B[7];
    assign stage0_r20_c6 = A[20] & B[6];
    assign stage0_r21_c5 = A[21] & B[5];
    assign stage0_r22_c4 = A[22] & B[4];
    assign stage0_r23_c3 = A[23] & B[3];
    assign stage0_r24_c2 = A[24] & B[2];
    assign stage0_r25_c1 = A[25] & B[1];
    assign stage0_r26_c0 = A[26] & B[0];
    assign stage0_r0_c27 = A[0] & B[27];
    assign stage0_r1_c26 = A[1] & B[26];
    assign stage0_r2_c25 = A[2] & B[25];
    assign stage0_r3_c24 = A[3] & B[24];
    assign stage0_r4_c23 = A[4] & B[23];
    assign stage0_r5_c22 = A[5] & B[22];
    assign stage0_r6_c21 = A[6] & B[21];
    assign stage0_r7_c20 = A[7] & B[20];
    assign stage0_r8_c19 = A[8] & B[19];
    assign stage0_r9_c18 = A[9] & B[18];
    assign stage0_r10_c17 = A[10] & B[17];
    assign stage0_r11_c16 = A[11] & B[16];
    assign stage0_r12_c15 = A[12] & B[15];
    assign stage0_r13_c14 = A[13] & B[14];
    assign stage0_r14_c13 = A[14] & B[13];
    assign stage0_r15_c12 = A[15] & B[12];
    assign stage0_r16_c11 = A[16] & B[11];
    assign stage0_r17_c10 = A[17] & B[10];
    assign stage0_r18_c9 = A[18] & B[9];
    assign stage0_r19_c8 = A[19] & B[8];
    assign stage0_r20_c7 = A[20] & B[7];
    assign stage0_r21_c6 = A[21] & B[6];
    assign stage0_r22_c5 = A[22] & B[5];
    assign stage0_r23_c4 = A[23] & B[4];
    assign stage0_r24_c3 = A[24] & B[3];
    assign stage0_r25_c2 = A[25] & B[2];
    assign stage0_r26_c1 = A[26] & B[1];
    assign stage0_r27_c0 = A[27] & B[0];
    assign stage0_r0_c28 = A[0] & B[28];
    assign stage0_r1_c27 = A[1] & B[27];
    assign stage0_r2_c26 = A[2] & B[26];
    assign stage0_r3_c25 = A[3] & B[25];
    assign stage0_r4_c24 = A[4] & B[24];
    assign stage0_r5_c23 = A[5] & B[23];
    assign stage0_r6_c22 = A[6] & B[22];
    assign stage0_r7_c21 = A[7] & B[21];
    assign stage0_r8_c20 = A[8] & B[20];
    assign stage0_r9_c19 = A[9] & B[19];
    assign stage0_r10_c18 = A[10] & B[18];
    assign stage0_r11_c17 = A[11] & B[17];
    assign stage0_r12_c16 = A[12] & B[16];
    assign stage0_r13_c15 = A[13] & B[15];
    assign stage0_r14_c14 = A[14] & B[14];
    assign stage0_r15_c13 = A[15] & B[13];
    assign stage0_r16_c12 = A[16] & B[12];
    assign stage0_r17_c11 = A[17] & B[11];
    assign stage0_r18_c10 = A[18] & B[10];
    assign stage0_r19_c9 = A[19] & B[9];
    assign stage0_r20_c8 = A[20] & B[8];
    assign stage0_r21_c7 = A[21] & B[7];
    assign stage0_r22_c6 = A[22] & B[6];
    assign stage0_r23_c5 = A[23] & B[5];
    assign stage0_r24_c4 = A[24] & B[4];
    assign stage0_r25_c3 = A[25] & B[3];
    assign stage0_r26_c2 = A[26] & B[2];
    assign stage0_r27_c1 = A[27] & B[1];
    assign stage0_r28_c0 = A[28] & B[0];
    assign stage0_r0_c29 = A[0] & B[29];
    assign stage0_r1_c28 = A[1] & B[28];
    assign stage0_r2_c27 = A[2] & B[27];
    assign stage0_r3_c26 = A[3] & B[26];
    assign stage0_r4_c25 = A[4] & B[25];
    assign stage0_r5_c24 = A[5] & B[24];
    assign stage0_r6_c23 = A[6] & B[23];
    assign stage0_r7_c22 = A[7] & B[22];
    assign stage0_r8_c21 = A[8] & B[21];
    assign stage0_r9_c20 = A[9] & B[20];
    assign stage0_r10_c19 = A[10] & B[19];
    assign stage0_r11_c18 = A[11] & B[18];
    assign stage0_r12_c17 = A[12] & B[17];
    assign stage0_r13_c16 = A[13] & B[16];
    assign stage0_r14_c15 = A[14] & B[15];
    assign stage0_r15_c14 = A[15] & B[14];
    assign stage0_r16_c13 = A[16] & B[13];
    assign stage0_r17_c12 = A[17] & B[12];
    assign stage0_r18_c11 = A[18] & B[11];
    assign stage0_r19_c10 = A[19] & B[10];
    assign stage0_r20_c9 = A[20] & B[9];
    assign stage0_r21_c8 = A[21] & B[8];
    assign stage0_r22_c7 = A[22] & B[7];
    assign stage0_r23_c6 = A[23] & B[6];
    assign stage0_r24_c5 = A[24] & B[5];
    assign stage0_r25_c4 = A[25] & B[4];
    assign stage0_r26_c3 = A[26] & B[3];
    assign stage0_r27_c2 = A[27] & B[2];
    assign stage0_r28_c1 = A[28] & B[1];
    assign stage0_r29_c0 = A[29] & B[0];
    assign stage0_r0_c30 = A[0] & B[30];
    assign stage0_r1_c29 = A[1] & B[29];
    assign stage0_r2_c28 = A[2] & B[28];
    assign stage0_r3_c27 = A[3] & B[27];
    assign stage0_r4_c26 = A[4] & B[26];
    assign stage0_r5_c25 = A[5] & B[25];
    assign stage0_r6_c24 = A[6] & B[24];
    assign stage0_r7_c23 = A[7] & B[23];
    assign stage0_r8_c22 = A[8] & B[22];
    assign stage0_r9_c21 = A[9] & B[21];
    assign stage0_r10_c20 = A[10] & B[20];
    assign stage0_r11_c19 = A[11] & B[19];
    assign stage0_r12_c18 = A[12] & B[18];
    assign stage0_r13_c17 = A[13] & B[17];
    assign stage0_r14_c16 = A[14] & B[16];
    assign stage0_r15_c15 = A[15] & B[15];
    assign stage0_r16_c14 = A[16] & B[14];
    assign stage0_r17_c13 = A[17] & B[13];
    assign stage0_r18_c12 = A[18] & B[12];
    assign stage0_r19_c11 = A[19] & B[11];
    assign stage0_r20_c10 = A[20] & B[10];
    assign stage0_r21_c9 = A[21] & B[9];
    assign stage0_r22_c8 = A[22] & B[8];
    assign stage0_r23_c7 = A[23] & B[7];
    assign stage0_r24_c6 = A[24] & B[6];
    assign stage0_r25_c5 = A[25] & B[5];
    assign stage0_r26_c4 = A[26] & B[4];
    assign stage0_r27_c3 = A[27] & B[3];
    assign stage0_r28_c2 = A[28] & B[2];
    assign stage0_r29_c1 = A[29] & B[1];
    assign stage0_r30_c0 = A[30] & B[0];
    assign stage0_r0_c31 = A[0] & B[31];
    assign stage0_r1_c30 = A[1] & B[30];
    assign stage0_r2_c29 = A[2] & B[29];
    assign stage0_r3_c28 = A[3] & B[28];
    assign stage0_r4_c27 = A[4] & B[27];
    assign stage0_r5_c26 = A[5] & B[26];
    assign stage0_r6_c25 = A[6] & B[25];
    assign stage0_r7_c24 = A[7] & B[24];
    assign stage0_r8_c23 = A[8] & B[23];
    assign stage0_r9_c22 = A[9] & B[22];
    assign stage0_r10_c21 = A[10] & B[21];
    assign stage0_r11_c20 = A[11] & B[20];
    assign stage0_r12_c19 = A[12] & B[19];
    assign stage0_r13_c18 = A[13] & B[18];
    assign stage0_r14_c17 = A[14] & B[17];
    assign stage0_r15_c16 = A[15] & B[16];
    assign stage0_r16_c15 = A[16] & B[15];
    assign stage0_r17_c14 = A[17] & B[14];
    assign stage0_r18_c13 = A[18] & B[13];
    assign stage0_r19_c12 = A[19] & B[12];
    assign stage0_r20_c11 = A[20] & B[11];
    assign stage0_r21_c10 = A[21] & B[10];
    assign stage0_r22_c9 = A[22] & B[9];
    assign stage0_r23_c8 = A[23] & B[8];
    assign stage0_r24_c7 = A[24] & B[7];
    assign stage0_r25_c6 = A[25] & B[6];
    assign stage0_r26_c5 = A[26] & B[5];
    assign stage0_r27_c4 = A[27] & B[4];
    assign stage0_r28_c3 = A[28] & B[3];
    assign stage0_r29_c2 = A[29] & B[2];
    assign stage0_r30_c1 = A[30] & B[1];
    assign stage0_r31_c0 = A[31] & B[0];
    assign stage0_r0_c32 = A[0] & B[32];
    assign stage0_r1_c31 = A[1] & B[31];
    assign stage0_r2_c30 = A[2] & B[30];
    assign stage0_r3_c29 = A[3] & B[29];
    assign stage0_r4_c28 = A[4] & B[28];
    assign stage0_r5_c27 = A[5] & B[27];
    assign stage0_r6_c26 = A[6] & B[26];
    assign stage0_r7_c25 = A[7] & B[25];
    assign stage0_r8_c24 = A[8] & B[24];
    assign stage0_r9_c23 = A[9] & B[23];
    assign stage0_r10_c22 = A[10] & B[22];
    assign stage0_r11_c21 = A[11] & B[21];
    assign stage0_r12_c20 = A[12] & B[20];
    assign stage0_r13_c19 = A[13] & B[19];
    assign stage0_r14_c18 = A[14] & B[18];
    assign stage0_r15_c17 = A[15] & B[17];
    assign stage0_r16_c16 = A[16] & B[16];
    assign stage0_r17_c15 = A[17] & B[15];
    assign stage0_r18_c14 = A[18] & B[14];
    assign stage0_r19_c13 = A[19] & B[13];
    assign stage0_r20_c12 = A[20] & B[12];
    assign stage0_r21_c11 = A[21] & B[11];
    assign stage0_r22_c10 = A[22] & B[10];
    assign stage0_r23_c9 = A[23] & B[9];
    assign stage0_r24_c8 = A[24] & B[8];
    assign stage0_r25_c7 = A[25] & B[7];
    assign stage0_r26_c6 = A[26] & B[6];
    assign stage0_r27_c5 = A[27] & B[5];
    assign stage0_r28_c4 = A[28] & B[4];
    assign stage0_r29_c3 = A[29] & B[3];
    assign stage0_r30_c2 = A[30] & B[2];
    assign stage0_r31_c1 = A[31] & B[1];
    assign stage0_r32_c0 = A[32] & B[0];
    assign stage0_r0_c33 = A[0] & B[33];
    assign stage0_r1_c32 = A[1] & B[32];
    assign stage0_r2_c31 = A[2] & B[31];
    assign stage0_r3_c30 = A[3] & B[30];
    assign stage0_r4_c29 = A[4] & B[29];
    assign stage0_r5_c28 = A[5] & B[28];
    assign stage0_r6_c27 = A[6] & B[27];
    assign stage0_r7_c26 = A[7] & B[26];
    assign stage0_r8_c25 = A[8] & B[25];
    assign stage0_r9_c24 = A[9] & B[24];
    assign stage0_r10_c23 = A[10] & B[23];
    assign stage0_r11_c22 = A[11] & B[22];
    assign stage0_r12_c21 = A[12] & B[21];
    assign stage0_r13_c20 = A[13] & B[20];
    assign stage0_r14_c19 = A[14] & B[19];
    assign stage0_r15_c18 = A[15] & B[18];
    assign stage0_r16_c17 = A[16] & B[17];
    assign stage0_r17_c16 = A[17] & B[16];
    assign stage0_r18_c15 = A[18] & B[15];
    assign stage0_r19_c14 = A[19] & B[14];
    assign stage0_r20_c13 = A[20] & B[13];
    assign stage0_r21_c12 = A[21] & B[12];
    assign stage0_r22_c11 = A[22] & B[11];
    assign stage0_r23_c10 = A[23] & B[10];
    assign stage0_r24_c9 = A[24] & B[9];
    assign stage0_r25_c8 = A[25] & B[8];
    assign stage0_r26_c7 = A[26] & B[7];
    assign stage0_r27_c6 = A[27] & B[6];
    assign stage0_r28_c5 = A[28] & B[5];
    assign stage0_r29_c4 = A[29] & B[4];
    assign stage0_r30_c3 = A[30] & B[3];
    assign stage0_r31_c2 = A[31] & B[2];
    assign stage0_r32_c1 = A[32] & B[1];
    assign stage0_r33_c0 = A[33] & B[0];
    assign stage0_r0_c34 = A[0] & B[34];
    assign stage0_r1_c33 = A[1] & B[33];
    assign stage0_r2_c32 = A[2] & B[32];
    assign stage0_r3_c31 = A[3] & B[31];
    assign stage0_r4_c30 = A[4] & B[30];
    assign stage0_r5_c29 = A[5] & B[29];
    assign stage0_r6_c28 = A[6] & B[28];
    assign stage0_r7_c27 = A[7] & B[27];
    assign stage0_r8_c26 = A[8] & B[26];
    assign stage0_r9_c25 = A[9] & B[25];
    assign stage0_r10_c24 = A[10] & B[24];
    assign stage0_r11_c23 = A[11] & B[23];
    assign stage0_r12_c22 = A[12] & B[22];
    assign stage0_r13_c21 = A[13] & B[21];
    assign stage0_r14_c20 = A[14] & B[20];
    assign stage0_r15_c19 = A[15] & B[19];
    assign stage0_r16_c18 = A[16] & B[18];
    assign stage0_r17_c17 = A[17] & B[17];
    assign stage0_r18_c16 = A[18] & B[16];
    assign stage0_r19_c15 = A[19] & B[15];
    assign stage0_r20_c14 = A[20] & B[14];
    assign stage0_r21_c13 = A[21] & B[13];
    assign stage0_r22_c12 = A[22] & B[12];
    assign stage0_r23_c11 = A[23] & B[11];
    assign stage0_r24_c10 = A[24] & B[10];
    assign stage0_r25_c9 = A[25] & B[9];
    assign stage0_r26_c8 = A[26] & B[8];
    assign stage0_r27_c7 = A[27] & B[7];
    assign stage0_r28_c6 = A[28] & B[6];
    assign stage0_r29_c5 = A[29] & B[5];
    assign stage0_r30_c4 = A[30] & B[4];
    assign stage0_r31_c3 = A[31] & B[3];
    assign stage0_r32_c2 = A[32] & B[2];
    assign stage0_r33_c1 = A[33] & B[1];
    assign stage0_r34_c0 = A[34] & B[0];
    assign stage0_r0_c35 = A[0] & B[35];
    assign stage0_r1_c34 = A[1] & B[34];
    assign stage0_r2_c33 = A[2] & B[33];
    assign stage0_r3_c32 = A[3] & B[32];
    assign stage0_r4_c31 = A[4] & B[31];
    assign stage0_r5_c30 = A[5] & B[30];
    assign stage0_r6_c29 = A[6] & B[29];
    assign stage0_r7_c28 = A[7] & B[28];
    assign stage0_r8_c27 = A[8] & B[27];
    assign stage0_r9_c26 = A[9] & B[26];
    assign stage0_r10_c25 = A[10] & B[25];
    assign stage0_r11_c24 = A[11] & B[24];
    assign stage0_r12_c23 = A[12] & B[23];
    assign stage0_r13_c22 = A[13] & B[22];
    assign stage0_r14_c21 = A[14] & B[21];
    assign stage0_r15_c20 = A[15] & B[20];
    assign stage0_r16_c19 = A[16] & B[19];
    assign stage0_r17_c18 = A[17] & B[18];
    assign stage0_r18_c17 = A[18] & B[17];
    assign stage0_r19_c16 = A[19] & B[16];
    assign stage0_r20_c15 = A[20] & B[15];
    assign stage0_r21_c14 = A[21] & B[14];
    assign stage0_r22_c13 = A[22] & B[13];
    assign stage0_r23_c12 = A[23] & B[12];
    assign stage0_r24_c11 = A[24] & B[11];
    assign stage0_r25_c10 = A[25] & B[10];
    assign stage0_r26_c9 = A[26] & B[9];
    assign stage0_r27_c8 = A[27] & B[8];
    assign stage0_r28_c7 = A[28] & B[7];
    assign stage0_r29_c6 = A[29] & B[6];
    assign stage0_r30_c5 = A[30] & B[5];
    assign stage0_r31_c4 = A[31] & B[4];
    assign stage0_r32_c3 = A[32] & B[3];
    assign stage0_r33_c2 = A[33] & B[2];
    assign stage0_r34_c1 = A[34] & B[1];
    assign stage0_r35_c0 = A[35] & B[0];
    assign stage0_r0_c36 = A[0] & B[36];
    assign stage0_r1_c35 = A[1] & B[35];
    assign stage0_r2_c34 = A[2] & B[34];
    assign stage0_r3_c33 = A[3] & B[33];
    assign stage0_r4_c32 = A[4] & B[32];
    assign stage0_r5_c31 = A[5] & B[31];
    assign stage0_r6_c30 = A[6] & B[30];
    assign stage0_r7_c29 = A[7] & B[29];
    assign stage0_r8_c28 = A[8] & B[28];
    assign stage0_r9_c27 = A[9] & B[27];
    assign stage0_r10_c26 = A[10] & B[26];
    assign stage0_r11_c25 = A[11] & B[25];
    assign stage0_r12_c24 = A[12] & B[24];
    assign stage0_r13_c23 = A[13] & B[23];
    assign stage0_r14_c22 = A[14] & B[22];
    assign stage0_r15_c21 = A[15] & B[21];
    assign stage0_r16_c20 = A[16] & B[20];
    assign stage0_r17_c19 = A[17] & B[19];
    assign stage0_r18_c18 = A[18] & B[18];
    assign stage0_r19_c17 = A[19] & B[17];
    assign stage0_r20_c16 = A[20] & B[16];
    assign stage0_r21_c15 = A[21] & B[15];
    assign stage0_r22_c14 = A[22] & B[14];
    assign stage0_r23_c13 = A[23] & B[13];
    assign stage0_r24_c12 = A[24] & B[12];
    assign stage0_r25_c11 = A[25] & B[11];
    assign stage0_r26_c10 = A[26] & B[10];
    assign stage0_r27_c9 = A[27] & B[9];
    assign stage0_r28_c8 = A[28] & B[8];
    assign stage0_r29_c7 = A[29] & B[7];
    assign stage0_r30_c6 = A[30] & B[6];
    assign stage0_r31_c5 = A[31] & B[5];
    assign stage0_r32_c4 = A[32] & B[4];
    assign stage0_r33_c3 = A[33] & B[3];
    assign stage0_r34_c2 = A[34] & B[2];
    assign stage0_r35_c1 = A[35] & B[1];
    assign stage0_r36_c0 = A[36] & B[0];
    assign stage0_r0_c37 = A[0] & B[37];
    assign stage0_r1_c36 = A[1] & B[36];
    assign stage0_r2_c35 = A[2] & B[35];
    assign stage0_r3_c34 = A[3] & B[34];
    assign stage0_r4_c33 = A[4] & B[33];
    assign stage0_r5_c32 = A[5] & B[32];
    assign stage0_r6_c31 = A[6] & B[31];
    assign stage0_r7_c30 = A[7] & B[30];
    assign stage0_r8_c29 = A[8] & B[29];
    assign stage0_r9_c28 = A[9] & B[28];
    assign stage0_r10_c27 = A[10] & B[27];
    assign stage0_r11_c26 = A[11] & B[26];
    assign stage0_r12_c25 = A[12] & B[25];
    assign stage0_r13_c24 = A[13] & B[24];
    assign stage0_r14_c23 = A[14] & B[23];
    assign stage0_r15_c22 = A[15] & B[22];
    assign stage0_r16_c21 = A[16] & B[21];
    assign stage0_r17_c20 = A[17] & B[20];
    assign stage0_r18_c19 = A[18] & B[19];
    assign stage0_r19_c18 = A[19] & B[18];
    assign stage0_r20_c17 = A[20] & B[17];
    assign stage0_r21_c16 = A[21] & B[16];
    assign stage0_r22_c15 = A[22] & B[15];
    assign stage0_r23_c14 = A[23] & B[14];
    assign stage0_r24_c13 = A[24] & B[13];
    assign stage0_r25_c12 = A[25] & B[12];
    assign stage0_r26_c11 = A[26] & B[11];
    assign stage0_r27_c10 = A[27] & B[10];
    assign stage0_r28_c9 = A[28] & B[9];
    assign stage0_r29_c8 = A[29] & B[8];
    assign stage0_r30_c7 = A[30] & B[7];
    assign stage0_r31_c6 = A[31] & B[6];
    assign stage0_r32_c5 = A[32] & B[5];
    assign stage0_r33_c4 = A[33] & B[4];
    assign stage0_r34_c3 = A[34] & B[3];
    assign stage0_r35_c2 = A[35] & B[2];
    assign stage0_r36_c1 = A[36] & B[1];
    assign stage0_r37_c0 = A[37] & B[0];
    assign stage0_r0_c38 = A[0] & B[38];
    assign stage0_r1_c37 = A[1] & B[37];
    assign stage0_r2_c36 = A[2] & B[36];
    assign stage0_r3_c35 = A[3] & B[35];
    assign stage0_r4_c34 = A[4] & B[34];
    assign stage0_r5_c33 = A[5] & B[33];
    assign stage0_r6_c32 = A[6] & B[32];
    assign stage0_r7_c31 = A[7] & B[31];
    assign stage0_r8_c30 = A[8] & B[30];
    assign stage0_r9_c29 = A[9] & B[29];
    assign stage0_r10_c28 = A[10] & B[28];
    assign stage0_r11_c27 = A[11] & B[27];
    assign stage0_r12_c26 = A[12] & B[26];
    assign stage0_r13_c25 = A[13] & B[25];
    assign stage0_r14_c24 = A[14] & B[24];
    assign stage0_r15_c23 = A[15] & B[23];
    assign stage0_r16_c22 = A[16] & B[22];
    assign stage0_r17_c21 = A[17] & B[21];
    assign stage0_r18_c20 = A[18] & B[20];
    assign stage0_r19_c19 = A[19] & B[19];
    assign stage0_r20_c18 = A[20] & B[18];
    assign stage0_r21_c17 = A[21] & B[17];
    assign stage0_r22_c16 = A[22] & B[16];
    assign stage0_r23_c15 = A[23] & B[15];
    assign stage0_r24_c14 = A[24] & B[14];
    assign stage0_r25_c13 = A[25] & B[13];
    assign stage0_r26_c12 = A[26] & B[12];
    assign stage0_r27_c11 = A[27] & B[11];
    assign stage0_r28_c10 = A[28] & B[10];
    assign stage0_r29_c9 = A[29] & B[9];
    assign stage0_r30_c8 = A[30] & B[8];
    assign stage0_r31_c7 = A[31] & B[7];
    assign stage0_r32_c6 = A[32] & B[6];
    assign stage0_r33_c5 = A[33] & B[5];
    assign stage0_r34_c4 = A[34] & B[4];
    assign stage0_r35_c3 = A[35] & B[3];
    assign stage0_r36_c2 = A[36] & B[2];
    assign stage0_r37_c1 = A[37] & B[1];
    assign stage0_r38_c0 = A[38] & B[0];
    assign stage0_r0_c39 = A[0] & B[39];
    assign stage0_r1_c38 = A[1] & B[38];
    assign stage0_r2_c37 = A[2] & B[37];
    assign stage0_r3_c36 = A[3] & B[36];
    assign stage0_r4_c35 = A[4] & B[35];
    assign stage0_r5_c34 = A[5] & B[34];
    assign stage0_r6_c33 = A[6] & B[33];
    assign stage0_r7_c32 = A[7] & B[32];
    assign stage0_r8_c31 = A[8] & B[31];
    assign stage0_r9_c30 = A[9] & B[30];
    assign stage0_r10_c29 = A[10] & B[29];
    assign stage0_r11_c28 = A[11] & B[28];
    assign stage0_r12_c27 = A[12] & B[27];
    assign stage0_r13_c26 = A[13] & B[26];
    assign stage0_r14_c25 = A[14] & B[25];
    assign stage0_r15_c24 = A[15] & B[24];
    assign stage0_r16_c23 = A[16] & B[23];
    assign stage0_r17_c22 = A[17] & B[22];
    assign stage0_r18_c21 = A[18] & B[21];
    assign stage0_r19_c20 = A[19] & B[20];
    assign stage0_r20_c19 = A[20] & B[19];
    assign stage0_r21_c18 = A[21] & B[18];
    assign stage0_r22_c17 = A[22] & B[17];
    assign stage0_r23_c16 = A[23] & B[16];
    assign stage0_r24_c15 = A[24] & B[15];
    assign stage0_r25_c14 = A[25] & B[14];
    assign stage0_r26_c13 = A[26] & B[13];
    assign stage0_r27_c12 = A[27] & B[12];
    assign stage0_r28_c11 = A[28] & B[11];
    assign stage0_r29_c10 = A[29] & B[10];
    assign stage0_r30_c9 = A[30] & B[9];
    assign stage0_r31_c8 = A[31] & B[8];
    assign stage0_r32_c7 = A[32] & B[7];
    assign stage0_r33_c6 = A[33] & B[6];
    assign stage0_r34_c5 = A[34] & B[5];
    assign stage0_r35_c4 = A[35] & B[4];
    assign stage0_r36_c3 = A[36] & B[3];
    assign stage0_r37_c2 = A[37] & B[2];
    assign stage0_r38_c1 = A[38] & B[1];
    assign stage0_r39_c0 = A[39] & B[0];
    assign stage0_r0_c40 = A[0] & B[40];
    assign stage0_r1_c39 = A[1] & B[39];
    assign stage0_r2_c38 = A[2] & B[38];
    assign stage0_r3_c37 = A[3] & B[37];
    assign stage0_r4_c36 = A[4] & B[36];
    assign stage0_r5_c35 = A[5] & B[35];
    assign stage0_r6_c34 = A[6] & B[34];
    assign stage0_r7_c33 = A[7] & B[33];
    assign stage0_r8_c32 = A[8] & B[32];
    assign stage0_r9_c31 = A[9] & B[31];
    assign stage0_r10_c30 = A[10] & B[30];
    assign stage0_r11_c29 = A[11] & B[29];
    assign stage0_r12_c28 = A[12] & B[28];
    assign stage0_r13_c27 = A[13] & B[27];
    assign stage0_r14_c26 = A[14] & B[26];
    assign stage0_r15_c25 = A[15] & B[25];
    assign stage0_r16_c24 = A[16] & B[24];
    assign stage0_r17_c23 = A[17] & B[23];
    assign stage0_r18_c22 = A[18] & B[22];
    assign stage0_r19_c21 = A[19] & B[21];
    assign stage0_r20_c20 = A[20] & B[20];
    assign stage0_r21_c19 = A[21] & B[19];
    assign stage0_r22_c18 = A[22] & B[18];
    assign stage0_r23_c17 = A[23] & B[17];
    assign stage0_r24_c16 = A[24] & B[16];
    assign stage0_r25_c15 = A[25] & B[15];
    assign stage0_r26_c14 = A[26] & B[14];
    assign stage0_r27_c13 = A[27] & B[13];
    assign stage0_r28_c12 = A[28] & B[12];
    assign stage0_r29_c11 = A[29] & B[11];
    assign stage0_r30_c10 = A[30] & B[10];
    assign stage0_r31_c9 = A[31] & B[9];
    assign stage0_r32_c8 = A[32] & B[8];
    assign stage0_r33_c7 = A[33] & B[7];
    assign stage0_r34_c6 = A[34] & B[6];
    assign stage0_r35_c5 = A[35] & B[5];
    assign stage0_r36_c4 = A[36] & B[4];
    assign stage0_r37_c3 = A[37] & B[3];
    assign stage0_r38_c2 = A[38] & B[2];
    assign stage0_r39_c1 = A[39] & B[1];
    assign stage0_r40_c0 = A[40] & B[0];
    assign stage0_r1_c40 = A[1] & B[40];
    assign stage0_r2_c39 = A[2] & B[39];
    assign stage0_r3_c38 = A[3] & B[38];
    assign stage0_r4_c37 = A[4] & B[37];
    assign stage0_r5_c36 = A[5] & B[36];
    assign stage0_r6_c35 = A[6] & B[35];
    assign stage0_r7_c34 = A[7] & B[34];
    assign stage0_r8_c33 = A[8] & B[33];
    assign stage0_r9_c32 = A[9] & B[32];
    assign stage0_r10_c31 = A[10] & B[31];
    assign stage0_r11_c30 = A[11] & B[30];
    assign stage0_r12_c29 = A[12] & B[29];
    assign stage0_r13_c28 = A[13] & B[28];
    assign stage0_r14_c27 = A[14] & B[27];
    assign stage0_r15_c26 = A[15] & B[26];
    assign stage0_r16_c25 = A[16] & B[25];
    assign stage0_r17_c24 = A[17] & B[24];
    assign stage0_r18_c23 = A[18] & B[23];
    assign stage0_r19_c22 = A[19] & B[22];
    assign stage0_r20_c21 = A[20] & B[21];
    assign stage0_r21_c20 = A[21] & B[20];
    assign stage0_r22_c19 = A[22] & B[19];
    assign stage0_r23_c18 = A[23] & B[18];
    assign stage0_r24_c17 = A[24] & B[17];
    assign stage0_r25_c16 = A[25] & B[16];
    assign stage0_r26_c15 = A[26] & B[15];
    assign stage0_r27_c14 = A[27] & B[14];
    assign stage0_r28_c13 = A[28] & B[13];
    assign stage0_r29_c12 = A[29] & B[12];
    assign stage0_r30_c11 = A[30] & B[11];
    assign stage0_r31_c10 = A[31] & B[10];
    assign stage0_r32_c9 = A[32] & B[9];
    assign stage0_r33_c8 = A[33] & B[8];
    assign stage0_r34_c7 = A[34] & B[7];
    assign stage0_r35_c6 = A[35] & B[6];
    assign stage0_r36_c5 = A[36] & B[5];
    assign stage0_r37_c4 = A[37] & B[4];
    assign stage0_r38_c3 = A[38] & B[3];
    assign stage0_r39_c2 = A[39] & B[2];
    assign stage0_r40_c1 = A[40] & B[1];
    assign stage0_r41_c0 = A[41] & B[0];
    assign stage0_r2_c40 = A[2] & B[40];
    assign stage0_r3_c39 = A[3] & B[39];
    assign stage0_r4_c38 = A[4] & B[38];
    assign stage0_r5_c37 = A[5] & B[37];
    assign stage0_r6_c36 = A[6] & B[36];
    assign stage0_r7_c35 = A[7] & B[35];
    assign stage0_r8_c34 = A[8] & B[34];
    assign stage0_r9_c33 = A[9] & B[33];
    assign stage0_r10_c32 = A[10] & B[32];
    assign stage0_r11_c31 = A[11] & B[31];
    assign stage0_r12_c30 = A[12] & B[30];
    assign stage0_r13_c29 = A[13] & B[29];
    assign stage0_r14_c28 = A[14] & B[28];
    assign stage0_r15_c27 = A[15] & B[27];
    assign stage0_r16_c26 = A[16] & B[26];
    assign stage0_r17_c25 = A[17] & B[25];
    assign stage0_r18_c24 = A[18] & B[24];
    assign stage0_r19_c23 = A[19] & B[23];
    assign stage0_r20_c22 = A[20] & B[22];
    assign stage0_r21_c21 = A[21] & B[21];
    assign stage0_r22_c20 = A[22] & B[20];
    assign stage0_r23_c19 = A[23] & B[19];
    assign stage0_r24_c18 = A[24] & B[18];
    assign stage0_r25_c17 = A[25] & B[17];
    assign stage0_r26_c16 = A[26] & B[16];
    assign stage0_r27_c15 = A[27] & B[15];
    assign stage0_r28_c14 = A[28] & B[14];
    assign stage0_r29_c13 = A[29] & B[13];
    assign stage0_r30_c12 = A[30] & B[12];
    assign stage0_r31_c11 = A[31] & B[11];
    assign stage0_r32_c10 = A[32] & B[10];
    assign stage0_r33_c9 = A[33] & B[9];
    assign stage0_r34_c8 = A[34] & B[8];
    assign stage0_r35_c7 = A[35] & B[7];
    assign stage0_r36_c6 = A[36] & B[6];
    assign stage0_r37_c5 = A[37] & B[5];
    assign stage0_r38_c4 = A[38] & B[4];
    assign stage0_r39_c3 = A[39] & B[3];
    assign stage0_r40_c2 = A[40] & B[2];
    assign stage0_r41_c1 = A[41] & B[1];
    assign stage0_r42_c0 = A[42] & B[0];
    assign stage0_r3_c40 = A[3] & B[40];
    assign stage0_r4_c39 = A[4] & B[39];
    assign stage0_r5_c38 = A[5] & B[38];
    assign stage0_r6_c37 = A[6] & B[37];
    assign stage0_r7_c36 = A[7] & B[36];
    assign stage0_r8_c35 = A[8] & B[35];
    assign stage0_r9_c34 = A[9] & B[34];
    assign stage0_r10_c33 = A[10] & B[33];
    assign stage0_r11_c32 = A[11] & B[32];
    assign stage0_r12_c31 = A[12] & B[31];
    assign stage0_r13_c30 = A[13] & B[30];
    assign stage0_r14_c29 = A[14] & B[29];
    assign stage0_r15_c28 = A[15] & B[28];
    assign stage0_r16_c27 = A[16] & B[27];
    assign stage0_r17_c26 = A[17] & B[26];
    assign stage0_r18_c25 = A[18] & B[25];
    assign stage0_r19_c24 = A[19] & B[24];
    assign stage0_r20_c23 = A[20] & B[23];
    assign stage0_r21_c22 = A[21] & B[22];
    assign stage0_r22_c21 = A[22] & B[21];
    assign stage0_r23_c20 = A[23] & B[20];
    assign stage0_r24_c19 = A[24] & B[19];
    assign stage0_r25_c18 = A[25] & B[18];
    assign stage0_r26_c17 = A[26] & B[17];
    assign stage0_r27_c16 = A[27] & B[16];
    assign stage0_r28_c15 = A[28] & B[15];
    assign stage0_r29_c14 = A[29] & B[14];
    assign stage0_r30_c13 = A[30] & B[13];
    assign stage0_r31_c12 = A[31] & B[12];
    assign stage0_r32_c11 = A[32] & B[11];
    assign stage0_r33_c10 = A[33] & B[10];
    assign stage0_r34_c9 = A[34] & B[9];
    assign stage0_r35_c8 = A[35] & B[8];
    assign stage0_r36_c7 = A[36] & B[7];
    assign stage0_r37_c6 = A[37] & B[6];
    assign stage0_r38_c5 = A[38] & B[5];
    assign stage0_r39_c4 = A[39] & B[4];
    assign stage0_r40_c3 = A[40] & B[3];
    assign stage0_r41_c2 = A[41] & B[2];
    assign stage0_r42_c1 = A[42] & B[1];
    assign stage0_r43_c0 = A[43] & B[0];
    assign stage0_r4_c40 = A[4] & B[40];
    assign stage0_r5_c39 = A[5] & B[39];
    assign stage0_r6_c38 = A[6] & B[38];
    assign stage0_r7_c37 = A[7] & B[37];
    assign stage0_r8_c36 = A[8] & B[36];
    assign stage0_r9_c35 = A[9] & B[35];
    assign stage0_r10_c34 = A[10] & B[34];
    assign stage0_r11_c33 = A[11] & B[33];
    assign stage0_r12_c32 = A[12] & B[32];
    assign stage0_r13_c31 = A[13] & B[31];
    assign stage0_r14_c30 = A[14] & B[30];
    assign stage0_r15_c29 = A[15] & B[29];
    assign stage0_r16_c28 = A[16] & B[28];
    assign stage0_r17_c27 = A[17] & B[27];
    assign stage0_r18_c26 = A[18] & B[26];
    assign stage0_r19_c25 = A[19] & B[25];
    assign stage0_r20_c24 = A[20] & B[24];
    assign stage0_r21_c23 = A[21] & B[23];
    assign stage0_r22_c22 = A[22] & B[22];
    assign stage0_r23_c21 = A[23] & B[21];
    assign stage0_r24_c20 = A[24] & B[20];
    assign stage0_r25_c19 = A[25] & B[19];
    assign stage0_r26_c18 = A[26] & B[18];
    assign stage0_r27_c17 = A[27] & B[17];
    assign stage0_r28_c16 = A[28] & B[16];
    assign stage0_r29_c15 = A[29] & B[15];
    assign stage0_r30_c14 = A[30] & B[14];
    assign stage0_r31_c13 = A[31] & B[13];
    assign stage0_r32_c12 = A[32] & B[12];
    assign stage0_r33_c11 = A[33] & B[11];
    assign stage0_r34_c10 = A[34] & B[10];
    assign stage0_r35_c9 = A[35] & B[9];
    assign stage0_r36_c8 = A[36] & B[8];
    assign stage0_r37_c7 = A[37] & B[7];
    assign stage0_r38_c6 = A[38] & B[6];
    assign stage0_r39_c5 = A[39] & B[5];
    assign stage0_r40_c4 = A[40] & B[4];
    assign stage0_r41_c3 = A[41] & B[3];
    assign stage0_r42_c2 = A[42] & B[2];
    assign stage0_r43_c1 = A[43] & B[1];
    assign stage0_r44_c0 = A[44] & B[0];
    assign stage0_r5_c40 = A[5] & B[40];
    assign stage0_r6_c39 = A[6] & B[39];
    assign stage0_r7_c38 = A[7] & B[38];
    assign stage0_r8_c37 = A[8] & B[37];
    assign stage0_r9_c36 = A[9] & B[36];
    assign stage0_r10_c35 = A[10] & B[35];
    assign stage0_r11_c34 = A[11] & B[34];
    assign stage0_r12_c33 = A[12] & B[33];
    assign stage0_r13_c32 = A[13] & B[32];
    assign stage0_r14_c31 = A[14] & B[31];
    assign stage0_r15_c30 = A[15] & B[30];
    assign stage0_r16_c29 = A[16] & B[29];
    assign stage0_r17_c28 = A[17] & B[28];
    assign stage0_r18_c27 = A[18] & B[27];
    assign stage0_r19_c26 = A[19] & B[26];
    assign stage0_r20_c25 = A[20] & B[25];
    assign stage0_r21_c24 = A[21] & B[24];
    assign stage0_r22_c23 = A[22] & B[23];
    assign stage0_r23_c22 = A[23] & B[22];
    assign stage0_r24_c21 = A[24] & B[21];
    assign stage0_r25_c20 = A[25] & B[20];
    assign stage0_r26_c19 = A[26] & B[19];
    assign stage0_r27_c18 = A[27] & B[18];
    assign stage0_r28_c17 = A[28] & B[17];
    assign stage0_r29_c16 = A[29] & B[16];
    assign stage0_r30_c15 = A[30] & B[15];
    assign stage0_r31_c14 = A[31] & B[14];
    assign stage0_r32_c13 = A[32] & B[13];
    assign stage0_r33_c12 = A[33] & B[12];
    assign stage0_r34_c11 = A[34] & B[11];
    assign stage0_r35_c10 = A[35] & B[10];
    assign stage0_r36_c9 = A[36] & B[9];
    assign stage0_r37_c8 = A[37] & B[8];
    assign stage0_r38_c7 = A[38] & B[7];
    assign stage0_r39_c6 = A[39] & B[6];
    assign stage0_r40_c5 = A[40] & B[5];
    assign stage0_r41_c4 = A[41] & B[4];
    assign stage0_r42_c3 = A[42] & B[3];
    assign stage0_r43_c2 = A[43] & B[2];
    assign stage0_r44_c1 = A[44] & B[1];
    assign stage0_r45_c0 = A[45] & B[0];
    assign stage0_r6_c40 = A[6] & B[40];
    assign stage0_r7_c39 = A[7] & B[39];
    assign stage0_r8_c38 = A[8] & B[38];
    assign stage0_r9_c37 = A[9] & B[37];
    assign stage0_r10_c36 = A[10] & B[36];
    assign stage0_r11_c35 = A[11] & B[35];
    assign stage0_r12_c34 = A[12] & B[34];
    assign stage0_r13_c33 = A[13] & B[33];
    assign stage0_r14_c32 = A[14] & B[32];
    assign stage0_r15_c31 = A[15] & B[31];
    assign stage0_r16_c30 = A[16] & B[30];
    assign stage0_r17_c29 = A[17] & B[29];
    assign stage0_r18_c28 = A[18] & B[28];
    assign stage0_r19_c27 = A[19] & B[27];
    assign stage0_r20_c26 = A[20] & B[26];
    assign stage0_r21_c25 = A[21] & B[25];
    assign stage0_r22_c24 = A[22] & B[24];
    assign stage0_r23_c23 = A[23] & B[23];
    assign stage0_r24_c22 = A[24] & B[22];
    assign stage0_r25_c21 = A[25] & B[21];
    assign stage0_r26_c20 = A[26] & B[20];
    assign stage0_r27_c19 = A[27] & B[19];
    assign stage0_r28_c18 = A[28] & B[18];
    assign stage0_r29_c17 = A[29] & B[17];
    assign stage0_r30_c16 = A[30] & B[16];
    assign stage0_r31_c15 = A[31] & B[15];
    assign stage0_r32_c14 = A[32] & B[14];
    assign stage0_r33_c13 = A[33] & B[13];
    assign stage0_r34_c12 = A[34] & B[12];
    assign stage0_r35_c11 = A[35] & B[11];
    assign stage0_r36_c10 = A[36] & B[10];
    assign stage0_r37_c9 = A[37] & B[9];
    assign stage0_r38_c8 = A[38] & B[8];
    assign stage0_r39_c7 = A[39] & B[7];
    assign stage0_r40_c6 = A[40] & B[6];
    assign stage0_r41_c5 = A[41] & B[5];
    assign stage0_r42_c4 = A[42] & B[4];
    assign stage0_r43_c3 = A[43] & B[3];
    assign stage0_r44_c2 = A[44] & B[2];
    assign stage0_r45_c1 = A[45] & B[1];
    assign stage0_r46_c0 = A[46] & B[0];
    assign stage0_r7_c40 = A[7] & B[40];
    assign stage0_r8_c39 = A[8] & B[39];
    assign stage0_r9_c38 = A[9] & B[38];
    assign stage0_r10_c37 = A[10] & B[37];
    assign stage0_r11_c36 = A[11] & B[36];
    assign stage0_r12_c35 = A[12] & B[35];
    assign stage0_r13_c34 = A[13] & B[34];
    assign stage0_r14_c33 = A[14] & B[33];
    assign stage0_r15_c32 = A[15] & B[32];
    assign stage0_r16_c31 = A[16] & B[31];
    assign stage0_r17_c30 = A[17] & B[30];
    assign stage0_r18_c29 = A[18] & B[29];
    assign stage0_r19_c28 = A[19] & B[28];
    assign stage0_r20_c27 = A[20] & B[27];
    assign stage0_r21_c26 = A[21] & B[26];
    assign stage0_r22_c25 = A[22] & B[25];
    assign stage0_r23_c24 = A[23] & B[24];
    assign stage0_r24_c23 = A[24] & B[23];
    assign stage0_r25_c22 = A[25] & B[22];
    assign stage0_r26_c21 = A[26] & B[21];
    assign stage0_r27_c20 = A[27] & B[20];
    assign stage0_r28_c19 = A[28] & B[19];
    assign stage0_r29_c18 = A[29] & B[18];
    assign stage0_r30_c17 = A[30] & B[17];
    assign stage0_r31_c16 = A[31] & B[16];
    assign stage0_r32_c15 = A[32] & B[15];
    assign stage0_r33_c14 = A[33] & B[14];
    assign stage0_r34_c13 = A[34] & B[13];
    assign stage0_r35_c12 = A[35] & B[12];
    assign stage0_r36_c11 = A[36] & B[11];
    assign stage0_r37_c10 = A[37] & B[10];
    assign stage0_r38_c9 = A[38] & B[9];
    assign stage0_r39_c8 = A[39] & B[8];
    assign stage0_r40_c7 = A[40] & B[7];
    assign stage0_r41_c6 = A[41] & B[6];
    assign stage0_r42_c5 = A[42] & B[5];
    assign stage0_r43_c4 = A[43] & B[4];
    assign stage0_r44_c3 = A[44] & B[3];
    assign stage0_r45_c2 = A[45] & B[2];
    assign stage0_r46_c1 = A[46] & B[1];
    assign stage0_r47_c0 = A[47] & B[0];
    assign stage0_r8_c40 = A[8] & B[40];
    assign stage0_r9_c39 = A[9] & B[39];
    assign stage0_r10_c38 = A[10] & B[38];
    assign stage0_r11_c37 = A[11] & B[37];
    assign stage0_r12_c36 = A[12] & B[36];
    assign stage0_r13_c35 = A[13] & B[35];
    assign stage0_r14_c34 = A[14] & B[34];
    assign stage0_r15_c33 = A[15] & B[33];
    assign stage0_r16_c32 = A[16] & B[32];
    assign stage0_r17_c31 = A[17] & B[31];
    assign stage0_r18_c30 = A[18] & B[30];
    assign stage0_r19_c29 = A[19] & B[29];
    assign stage0_r20_c28 = A[20] & B[28];
    assign stage0_r21_c27 = A[21] & B[27];
    assign stage0_r22_c26 = A[22] & B[26];
    assign stage0_r23_c25 = A[23] & B[25];
    assign stage0_r24_c24 = A[24] & B[24];
    assign stage0_r25_c23 = A[25] & B[23];
    assign stage0_r26_c22 = A[26] & B[22];
    assign stage0_r27_c21 = A[27] & B[21];
    assign stage0_r28_c20 = A[28] & B[20];
    assign stage0_r29_c19 = A[29] & B[19];
    assign stage0_r30_c18 = A[30] & B[18];
    assign stage0_r31_c17 = A[31] & B[17];
    assign stage0_r32_c16 = A[32] & B[16];
    assign stage0_r33_c15 = A[33] & B[15];
    assign stage0_r34_c14 = A[34] & B[14];
    assign stage0_r35_c13 = A[35] & B[13];
    assign stage0_r36_c12 = A[36] & B[12];
    assign stage0_r37_c11 = A[37] & B[11];
    assign stage0_r38_c10 = A[38] & B[10];
    assign stage0_r39_c9 = A[39] & B[9];
    assign stage0_r40_c8 = A[40] & B[8];
    assign stage0_r41_c7 = A[41] & B[7];
    assign stage0_r42_c6 = A[42] & B[6];
    assign stage0_r43_c5 = A[43] & B[5];
    assign stage0_r44_c4 = A[44] & B[4];
    assign stage0_r45_c3 = A[45] & B[3];
    assign stage0_r46_c2 = A[46] & B[2];
    assign stage0_r47_c1 = A[47] & B[1];
    assign stage0_r48_c0 = A[48] & B[0];
    assign stage0_r9_c40 = A[9] & B[40];
    assign stage0_r10_c39 = A[10] & B[39];
    assign stage0_r11_c38 = A[11] & B[38];
    assign stage0_r12_c37 = A[12] & B[37];
    assign stage0_r13_c36 = A[13] & B[36];
    assign stage0_r14_c35 = A[14] & B[35];
    assign stage0_r15_c34 = A[15] & B[34];
    assign stage0_r16_c33 = A[16] & B[33];
    assign stage0_r17_c32 = A[17] & B[32];
    assign stage0_r18_c31 = A[18] & B[31];
    assign stage0_r19_c30 = A[19] & B[30];
    assign stage0_r20_c29 = A[20] & B[29];
    assign stage0_r21_c28 = A[21] & B[28];
    assign stage0_r22_c27 = A[22] & B[27];
    assign stage0_r23_c26 = A[23] & B[26];
    assign stage0_r24_c25 = A[24] & B[25];
    assign stage0_r25_c24 = A[25] & B[24];
    assign stage0_r26_c23 = A[26] & B[23];
    assign stage0_r27_c22 = A[27] & B[22];
    assign stage0_r28_c21 = A[28] & B[21];
    assign stage0_r29_c20 = A[29] & B[20];
    assign stage0_r30_c19 = A[30] & B[19];
    assign stage0_r31_c18 = A[31] & B[18];
    assign stage0_r32_c17 = A[32] & B[17];
    assign stage0_r33_c16 = A[33] & B[16];
    assign stage0_r34_c15 = A[34] & B[15];
    assign stage0_r35_c14 = A[35] & B[14];
    assign stage0_r36_c13 = A[36] & B[13];
    assign stage0_r37_c12 = A[37] & B[12];
    assign stage0_r38_c11 = A[38] & B[11];
    assign stage0_r39_c10 = A[39] & B[10];
    assign stage0_r40_c9 = A[40] & B[9];
    assign stage0_r41_c8 = A[41] & B[8];
    assign stage0_r42_c7 = A[42] & B[7];
    assign stage0_r43_c6 = A[43] & B[6];
    assign stage0_r44_c5 = A[44] & B[5];
    assign stage0_r45_c4 = A[45] & B[4];
    assign stage0_r46_c3 = A[46] & B[3];
    assign stage0_r47_c2 = A[47] & B[2];
    assign stage0_r48_c1 = A[48] & B[1];
    assign stage0_r49_c0 = A[49] & B[0];
    assign stage0_r10_c40 = A[10] & B[40];
    assign stage0_r11_c39 = A[11] & B[39];
    assign stage0_r12_c38 = A[12] & B[38];
    assign stage0_r13_c37 = A[13] & B[37];
    assign stage0_r14_c36 = A[14] & B[36];
    assign stage0_r15_c35 = A[15] & B[35];
    assign stage0_r16_c34 = A[16] & B[34];
    assign stage0_r17_c33 = A[17] & B[33];
    assign stage0_r18_c32 = A[18] & B[32];
    assign stage0_r19_c31 = A[19] & B[31];
    assign stage0_r20_c30 = A[20] & B[30];
    assign stage0_r21_c29 = A[21] & B[29];
    assign stage0_r22_c28 = A[22] & B[28];
    assign stage0_r23_c27 = A[23] & B[27];
    assign stage0_r24_c26 = A[24] & B[26];
    assign stage0_r25_c25 = A[25] & B[25];
    assign stage0_r26_c24 = A[26] & B[24];
    assign stage0_r27_c23 = A[27] & B[23];
    assign stage0_r28_c22 = A[28] & B[22];
    assign stage0_r29_c21 = A[29] & B[21];
    assign stage0_r30_c20 = A[30] & B[20];
    assign stage0_r31_c19 = A[31] & B[19];
    assign stage0_r32_c18 = A[32] & B[18];
    assign stage0_r33_c17 = A[33] & B[17];
    assign stage0_r34_c16 = A[34] & B[16];
    assign stage0_r35_c15 = A[35] & B[15];
    assign stage0_r36_c14 = A[36] & B[14];
    assign stage0_r37_c13 = A[37] & B[13];
    assign stage0_r38_c12 = A[38] & B[12];
    assign stage0_r39_c11 = A[39] & B[11];
    assign stage0_r40_c10 = A[40] & B[10];
    assign stage0_r41_c9 = A[41] & B[9];
    assign stage0_r42_c8 = A[42] & B[8];
    assign stage0_r43_c7 = A[43] & B[7];
    assign stage0_r44_c6 = A[44] & B[6];
    assign stage0_r45_c5 = A[45] & B[5];
    assign stage0_r46_c4 = A[46] & B[4];
    assign stage0_r47_c3 = A[47] & B[3];
    assign stage0_r48_c2 = A[48] & B[2];
    assign stage0_r49_c1 = A[49] & B[1];
    assign stage0_r50_c0 = A[50] & B[0];
    assign stage0_r11_c40 = A[11] & B[40];
    assign stage0_r12_c39 = A[12] & B[39];
    assign stage0_r13_c38 = A[13] & B[38];
    assign stage0_r14_c37 = A[14] & B[37];
    assign stage0_r15_c36 = A[15] & B[36];
    assign stage0_r16_c35 = A[16] & B[35];
    assign stage0_r17_c34 = A[17] & B[34];
    assign stage0_r18_c33 = A[18] & B[33];
    assign stage0_r19_c32 = A[19] & B[32];
    assign stage0_r20_c31 = A[20] & B[31];
    assign stage0_r21_c30 = A[21] & B[30];
    assign stage0_r22_c29 = A[22] & B[29];
    assign stage0_r23_c28 = A[23] & B[28];
    assign stage0_r24_c27 = A[24] & B[27];
    assign stage0_r25_c26 = A[25] & B[26];
    assign stage0_r26_c25 = A[26] & B[25];
    assign stage0_r27_c24 = A[27] & B[24];
    assign stage0_r28_c23 = A[28] & B[23];
    assign stage0_r29_c22 = A[29] & B[22];
    assign stage0_r30_c21 = A[30] & B[21];
    assign stage0_r31_c20 = A[31] & B[20];
    assign stage0_r32_c19 = A[32] & B[19];
    assign stage0_r33_c18 = A[33] & B[18];
    assign stage0_r34_c17 = A[34] & B[17];
    assign stage0_r35_c16 = A[35] & B[16];
    assign stage0_r36_c15 = A[36] & B[15];
    assign stage0_r37_c14 = A[37] & B[14];
    assign stage0_r38_c13 = A[38] & B[13];
    assign stage0_r39_c12 = A[39] & B[12];
    assign stage0_r40_c11 = A[40] & B[11];
    assign stage0_r41_c10 = A[41] & B[10];
    assign stage0_r42_c9 = A[42] & B[9];
    assign stage0_r43_c8 = A[43] & B[8];
    assign stage0_r44_c7 = A[44] & B[7];
    assign stage0_r45_c6 = A[45] & B[6];
    assign stage0_r46_c5 = A[46] & B[5];
    assign stage0_r47_c4 = A[47] & B[4];
    assign stage0_r48_c3 = A[48] & B[3];
    assign stage0_r49_c2 = A[49] & B[2];
    assign stage0_r50_c1 = A[50] & B[1];
    assign stage0_r51_c0 = A[51] & B[0];
    assign stage0_r12_c40 = A[12] & B[40];
    assign stage0_r13_c39 = A[13] & B[39];
    assign stage0_r14_c38 = A[14] & B[38];
    assign stage0_r15_c37 = A[15] & B[37];
    assign stage0_r16_c36 = A[16] & B[36];
    assign stage0_r17_c35 = A[17] & B[35];
    assign stage0_r18_c34 = A[18] & B[34];
    assign stage0_r19_c33 = A[19] & B[33];
    assign stage0_r20_c32 = A[20] & B[32];
    assign stage0_r21_c31 = A[21] & B[31];
    assign stage0_r22_c30 = A[22] & B[30];
    assign stage0_r23_c29 = A[23] & B[29];
    assign stage0_r24_c28 = A[24] & B[28];
    assign stage0_r25_c27 = A[25] & B[27];
    assign stage0_r26_c26 = A[26] & B[26];
    assign stage0_r27_c25 = A[27] & B[25];
    assign stage0_r28_c24 = A[28] & B[24];
    assign stage0_r29_c23 = A[29] & B[23];
    assign stage0_r30_c22 = A[30] & B[22];
    assign stage0_r31_c21 = A[31] & B[21];
    assign stage0_r32_c20 = A[32] & B[20];
    assign stage0_r33_c19 = A[33] & B[19];
    assign stage0_r34_c18 = A[34] & B[18];
    assign stage0_r35_c17 = A[35] & B[17];
    assign stage0_r36_c16 = A[36] & B[16];
    assign stage0_r37_c15 = A[37] & B[15];
    assign stage0_r38_c14 = A[38] & B[14];
    assign stage0_r39_c13 = A[39] & B[13];
    assign stage0_r40_c12 = A[40] & B[12];
    assign stage0_r41_c11 = A[41] & B[11];
    assign stage0_r42_c10 = A[42] & B[10];
    assign stage0_r43_c9 = A[43] & B[9];
    assign stage0_r44_c8 = A[44] & B[8];
    assign stage0_r45_c7 = A[45] & B[7];
    assign stage0_r46_c6 = A[46] & B[6];
    assign stage0_r47_c5 = A[47] & B[5];
    assign stage0_r48_c4 = A[48] & B[4];
    assign stage0_r49_c3 = A[49] & B[3];
    assign stage0_r50_c2 = A[50] & B[2];
    assign stage0_r51_c1 = A[51] & B[1];
    assign stage0_r52_c0 = A[52] & B[0];
    assign stage0_r13_c40 = A[13] & B[40];
    assign stage0_r14_c39 = A[14] & B[39];
    assign stage0_r15_c38 = A[15] & B[38];
    assign stage0_r16_c37 = A[16] & B[37];
    assign stage0_r17_c36 = A[17] & B[36];
    assign stage0_r18_c35 = A[18] & B[35];
    assign stage0_r19_c34 = A[19] & B[34];
    assign stage0_r20_c33 = A[20] & B[33];
    assign stage0_r21_c32 = A[21] & B[32];
    assign stage0_r22_c31 = A[22] & B[31];
    assign stage0_r23_c30 = A[23] & B[30];
    assign stage0_r24_c29 = A[24] & B[29];
    assign stage0_r25_c28 = A[25] & B[28];
    assign stage0_r26_c27 = A[26] & B[27];
    assign stage0_r27_c26 = A[27] & B[26];
    assign stage0_r28_c25 = A[28] & B[25];
    assign stage0_r29_c24 = A[29] & B[24];
    assign stage0_r30_c23 = A[30] & B[23];
    assign stage0_r31_c22 = A[31] & B[22];
    assign stage0_r32_c21 = A[32] & B[21];
    assign stage0_r33_c20 = A[33] & B[20];
    assign stage0_r34_c19 = A[34] & B[19];
    assign stage0_r35_c18 = A[35] & B[18];
    assign stage0_r36_c17 = A[36] & B[17];
    assign stage0_r37_c16 = A[37] & B[16];
    assign stage0_r38_c15 = A[38] & B[15];
    assign stage0_r39_c14 = A[39] & B[14];
    assign stage0_r40_c13 = A[40] & B[13];
    assign stage0_r41_c12 = A[41] & B[12];
    assign stage0_r42_c11 = A[42] & B[11];
    assign stage0_r43_c10 = A[43] & B[10];
    assign stage0_r44_c9 = A[44] & B[9];
    assign stage0_r45_c8 = A[45] & B[8];
    assign stage0_r46_c7 = A[46] & B[7];
    assign stage0_r47_c6 = A[47] & B[6];
    assign stage0_r48_c5 = A[48] & B[5];
    assign stage0_r49_c4 = A[49] & B[4];
    assign stage0_r50_c3 = A[50] & B[3];
    assign stage0_r51_c2 = A[51] & B[2];
    assign stage0_r52_c1 = A[52] & B[1];
    assign stage0_r53_c0 = A[53] & B[0];
    assign stage0_r14_c40 = A[14] & B[40];
    assign stage0_r15_c39 = A[15] & B[39];
    assign stage0_r16_c38 = A[16] & B[38];
    assign stage0_r17_c37 = A[17] & B[37];
    assign stage0_r18_c36 = A[18] & B[36];
    assign stage0_r19_c35 = A[19] & B[35];
    assign stage0_r20_c34 = A[20] & B[34];
    assign stage0_r21_c33 = A[21] & B[33];
    assign stage0_r22_c32 = A[22] & B[32];
    assign stage0_r23_c31 = A[23] & B[31];
    assign stage0_r24_c30 = A[24] & B[30];
    assign stage0_r25_c29 = A[25] & B[29];
    assign stage0_r26_c28 = A[26] & B[28];
    assign stage0_r27_c27 = A[27] & B[27];
    assign stage0_r28_c26 = A[28] & B[26];
    assign stage0_r29_c25 = A[29] & B[25];
    assign stage0_r30_c24 = A[30] & B[24];
    assign stage0_r31_c23 = A[31] & B[23];
    assign stage0_r32_c22 = A[32] & B[22];
    assign stage0_r33_c21 = A[33] & B[21];
    assign stage0_r34_c20 = A[34] & B[20];
    assign stage0_r35_c19 = A[35] & B[19];
    assign stage0_r36_c18 = A[36] & B[18];
    assign stage0_r37_c17 = A[37] & B[17];
    assign stage0_r38_c16 = A[38] & B[16];
    assign stage0_r39_c15 = A[39] & B[15];
    assign stage0_r40_c14 = A[40] & B[14];
    assign stage0_r41_c13 = A[41] & B[13];
    assign stage0_r42_c12 = A[42] & B[12];
    assign stage0_r43_c11 = A[43] & B[11];
    assign stage0_r44_c10 = A[44] & B[10];
    assign stage0_r45_c9 = A[45] & B[9];
    assign stage0_r46_c8 = A[46] & B[8];
    assign stage0_r47_c7 = A[47] & B[7];
    assign stage0_r48_c6 = A[48] & B[6];
    assign stage0_r49_c5 = A[49] & B[5];
    assign stage0_r50_c4 = A[50] & B[4];
    assign stage0_r51_c3 = A[51] & B[3];
    assign stage0_r52_c2 = A[52] & B[2];
    assign stage0_r53_c1 = A[53] & B[1];
    assign stage0_r54_c0 = A[54] & B[0];
    assign stage0_r15_c40 = A[15] & B[40];
    assign stage0_r16_c39 = A[16] & B[39];
    assign stage0_r17_c38 = A[17] & B[38];
    assign stage0_r18_c37 = A[18] & B[37];
    assign stage0_r19_c36 = A[19] & B[36];
    assign stage0_r20_c35 = A[20] & B[35];
    assign stage0_r21_c34 = A[21] & B[34];
    assign stage0_r22_c33 = A[22] & B[33];
    assign stage0_r23_c32 = A[23] & B[32];
    assign stage0_r24_c31 = A[24] & B[31];
    assign stage0_r25_c30 = A[25] & B[30];
    assign stage0_r26_c29 = A[26] & B[29];
    assign stage0_r27_c28 = A[27] & B[28];
    assign stage0_r28_c27 = A[28] & B[27];
    assign stage0_r29_c26 = A[29] & B[26];
    assign stage0_r30_c25 = A[30] & B[25];
    assign stage0_r31_c24 = A[31] & B[24];
    assign stage0_r32_c23 = A[32] & B[23];
    assign stage0_r33_c22 = A[33] & B[22];
    assign stage0_r34_c21 = A[34] & B[21];
    assign stage0_r35_c20 = A[35] & B[20];
    assign stage0_r36_c19 = A[36] & B[19];
    assign stage0_r37_c18 = A[37] & B[18];
    assign stage0_r38_c17 = A[38] & B[17];
    assign stage0_r39_c16 = A[39] & B[16];
    assign stage0_r40_c15 = A[40] & B[15];
    assign stage0_r41_c14 = A[41] & B[14];
    assign stage0_r42_c13 = A[42] & B[13];
    assign stage0_r43_c12 = A[43] & B[12];
    assign stage0_r44_c11 = A[44] & B[11];
    assign stage0_r45_c10 = A[45] & B[10];
    assign stage0_r46_c9 = A[46] & B[9];
    assign stage0_r47_c8 = A[47] & B[8];
    assign stage0_r48_c7 = A[48] & B[7];
    assign stage0_r49_c6 = A[49] & B[6];
    assign stage0_r50_c5 = A[50] & B[5];
    assign stage0_r51_c4 = A[51] & B[4];
    assign stage0_r52_c3 = A[52] & B[3];
    assign stage0_r53_c2 = A[53] & B[2];
    assign stage0_r54_c1 = A[54] & B[1];
    assign stage0_r55_c0 = A[55] & B[0];
    assign stage0_r16_c40 = A[16] & B[40];
    assign stage0_r17_c39 = A[17] & B[39];
    assign stage0_r18_c38 = A[18] & B[38];
    assign stage0_r19_c37 = A[19] & B[37];
    assign stage0_r20_c36 = A[20] & B[36];
    assign stage0_r21_c35 = A[21] & B[35];
    assign stage0_r22_c34 = A[22] & B[34];
    assign stage0_r23_c33 = A[23] & B[33];
    assign stage0_r24_c32 = A[24] & B[32];
    assign stage0_r25_c31 = A[25] & B[31];
    assign stage0_r26_c30 = A[26] & B[30];
    assign stage0_r27_c29 = A[27] & B[29];
    assign stage0_r28_c28 = A[28] & B[28];
    assign stage0_r29_c27 = A[29] & B[27];
    assign stage0_r30_c26 = A[30] & B[26];
    assign stage0_r31_c25 = A[31] & B[25];
    assign stage0_r32_c24 = A[32] & B[24];
    assign stage0_r33_c23 = A[33] & B[23];
    assign stage0_r34_c22 = A[34] & B[22];
    assign stage0_r35_c21 = A[35] & B[21];
    assign stage0_r36_c20 = A[36] & B[20];
    assign stage0_r37_c19 = A[37] & B[19];
    assign stage0_r38_c18 = A[38] & B[18];
    assign stage0_r39_c17 = A[39] & B[17];
    assign stage0_r40_c16 = A[40] & B[16];
    assign stage0_r41_c15 = A[41] & B[15];
    assign stage0_r42_c14 = A[42] & B[14];
    assign stage0_r43_c13 = A[43] & B[13];
    assign stage0_r44_c12 = A[44] & B[12];
    assign stage0_r45_c11 = A[45] & B[11];
    assign stage0_r46_c10 = A[46] & B[10];
    assign stage0_r47_c9 = A[47] & B[9];
    assign stage0_r48_c8 = A[48] & B[8];
    assign stage0_r49_c7 = A[49] & B[7];
    assign stage0_r50_c6 = A[50] & B[6];
    assign stage0_r51_c5 = A[51] & B[5];
    assign stage0_r52_c4 = A[52] & B[4];
    assign stage0_r53_c3 = A[53] & B[3];
    assign stage0_r54_c2 = A[54] & B[2];
    assign stage0_r55_c1 = A[55] & B[1];
    assign stage0_r56_c0 = A[56] & B[0];
    assign stage0_r17_c40 = A[17] & B[40];
    assign stage0_r18_c39 = A[18] & B[39];
    assign stage0_r19_c38 = A[19] & B[38];
    assign stage0_r20_c37 = A[20] & B[37];
    assign stage0_r21_c36 = A[21] & B[36];
    assign stage0_r22_c35 = A[22] & B[35];
    assign stage0_r23_c34 = A[23] & B[34];
    assign stage0_r24_c33 = A[24] & B[33];
    assign stage0_r25_c32 = A[25] & B[32];
    assign stage0_r26_c31 = A[26] & B[31];
    assign stage0_r27_c30 = A[27] & B[30];
    assign stage0_r28_c29 = A[28] & B[29];
    assign stage0_r29_c28 = A[29] & B[28];
    assign stage0_r30_c27 = A[30] & B[27];
    assign stage0_r31_c26 = A[31] & B[26];
    assign stage0_r32_c25 = A[32] & B[25];
    assign stage0_r33_c24 = A[33] & B[24];
    assign stage0_r34_c23 = A[34] & B[23];
    assign stage0_r35_c22 = A[35] & B[22];
    assign stage0_r36_c21 = A[36] & B[21];
    assign stage0_r37_c20 = A[37] & B[20];
    assign stage0_r38_c19 = A[38] & B[19];
    assign stage0_r39_c18 = A[39] & B[18];
    assign stage0_r40_c17 = A[40] & B[17];
    assign stage0_r41_c16 = A[41] & B[16];
    assign stage0_r42_c15 = A[42] & B[15];
    assign stage0_r43_c14 = A[43] & B[14];
    assign stage0_r44_c13 = A[44] & B[13];
    assign stage0_r45_c12 = A[45] & B[12];
    assign stage0_r46_c11 = A[46] & B[11];
    assign stage0_r47_c10 = A[47] & B[10];
    assign stage0_r48_c9 = A[48] & B[9];
    assign stage0_r49_c8 = A[49] & B[8];
    assign stage0_r50_c7 = A[50] & B[7];
    assign stage0_r51_c6 = A[51] & B[6];
    assign stage0_r52_c5 = A[52] & B[5];
    assign stage0_r53_c4 = A[53] & B[4];
    assign stage0_r54_c3 = A[54] & B[3];
    assign stage0_r55_c2 = A[55] & B[2];
    assign stage0_r56_c1 = A[56] & B[1];
    assign stage0_r57_c0 = A[57] & B[0];
    assign stage0_r18_c40 = A[18] & B[40];
    assign stage0_r19_c39 = A[19] & B[39];
    assign stage0_r20_c38 = A[20] & B[38];
    assign stage0_r21_c37 = A[21] & B[37];
    assign stage0_r22_c36 = A[22] & B[36];
    assign stage0_r23_c35 = A[23] & B[35];
    assign stage0_r24_c34 = A[24] & B[34];
    assign stage0_r25_c33 = A[25] & B[33];
    assign stage0_r26_c32 = A[26] & B[32];
    assign stage0_r27_c31 = A[27] & B[31];
    assign stage0_r28_c30 = A[28] & B[30];
    assign stage0_r29_c29 = A[29] & B[29];
    assign stage0_r30_c28 = A[30] & B[28];
    assign stage0_r31_c27 = A[31] & B[27];
    assign stage0_r32_c26 = A[32] & B[26];
    assign stage0_r33_c25 = A[33] & B[25];
    assign stage0_r34_c24 = A[34] & B[24];
    assign stage0_r35_c23 = A[35] & B[23];
    assign stage0_r36_c22 = A[36] & B[22];
    assign stage0_r37_c21 = A[37] & B[21];
    assign stage0_r38_c20 = A[38] & B[20];
    assign stage0_r39_c19 = A[39] & B[19];
    assign stage0_r40_c18 = A[40] & B[18];
    assign stage0_r41_c17 = A[41] & B[17];
    assign stage0_r42_c16 = A[42] & B[16];
    assign stage0_r43_c15 = A[43] & B[15];
    assign stage0_r44_c14 = A[44] & B[14];
    assign stage0_r45_c13 = A[45] & B[13];
    assign stage0_r46_c12 = A[46] & B[12];
    assign stage0_r47_c11 = A[47] & B[11];
    assign stage0_r48_c10 = A[48] & B[10];
    assign stage0_r49_c9 = A[49] & B[9];
    assign stage0_r50_c8 = A[50] & B[8];
    assign stage0_r51_c7 = A[51] & B[7];
    assign stage0_r52_c6 = A[52] & B[6];
    assign stage0_r53_c5 = A[53] & B[5];
    assign stage0_r54_c4 = A[54] & B[4];
    assign stage0_r55_c3 = A[55] & B[3];
    assign stage0_r56_c2 = A[56] & B[2];
    assign stage0_r57_c1 = A[57] & B[1];
    assign stage0_r58_c0 = A[58] & B[0];
    assign stage0_r19_c40 = A[19] & B[40];
    assign stage0_r20_c39 = A[20] & B[39];
    assign stage0_r21_c38 = A[21] & B[38];
    assign stage0_r22_c37 = A[22] & B[37];
    assign stage0_r23_c36 = A[23] & B[36];
    assign stage0_r24_c35 = A[24] & B[35];
    assign stage0_r25_c34 = A[25] & B[34];
    assign stage0_r26_c33 = A[26] & B[33];
    assign stage0_r27_c32 = A[27] & B[32];
    assign stage0_r28_c31 = A[28] & B[31];
    assign stage0_r29_c30 = A[29] & B[30];
    assign stage0_r30_c29 = A[30] & B[29];
    assign stage0_r31_c28 = A[31] & B[28];
    assign stage0_r32_c27 = A[32] & B[27];
    assign stage0_r33_c26 = A[33] & B[26];
    assign stage0_r34_c25 = A[34] & B[25];
    assign stage0_r35_c24 = A[35] & B[24];
    assign stage0_r36_c23 = A[36] & B[23];
    assign stage0_r37_c22 = A[37] & B[22];
    assign stage0_r38_c21 = A[38] & B[21];
    assign stage0_r39_c20 = A[39] & B[20];
    assign stage0_r40_c19 = A[40] & B[19];
    assign stage0_r41_c18 = A[41] & B[18];
    assign stage0_r42_c17 = A[42] & B[17];
    assign stage0_r43_c16 = A[43] & B[16];
    assign stage0_r44_c15 = A[44] & B[15];
    assign stage0_r45_c14 = A[45] & B[14];
    assign stage0_r46_c13 = A[46] & B[13];
    assign stage0_r47_c12 = A[47] & B[12];
    assign stage0_r48_c11 = A[48] & B[11];
    assign stage0_r49_c10 = A[49] & B[10];
    assign stage0_r50_c9 = A[50] & B[9];
    assign stage0_r51_c8 = A[51] & B[8];
    assign stage0_r52_c7 = A[52] & B[7];
    assign stage0_r53_c6 = A[53] & B[6];
    assign stage0_r54_c5 = A[54] & B[5];
    assign stage0_r55_c4 = A[55] & B[4];
    assign stage0_r56_c3 = A[56] & B[3];
    assign stage0_r57_c2 = A[57] & B[2];
    assign stage0_r58_c1 = A[58] & B[1];
    assign stage0_r59_c0 = A[59] & B[0];
    assign stage0_r20_c40 = A[20] & B[40];
    assign stage0_r21_c39 = A[21] & B[39];
    assign stage0_r22_c38 = A[22] & B[38];
    assign stage0_r23_c37 = A[23] & B[37];
    assign stage0_r24_c36 = A[24] & B[36];
    assign stage0_r25_c35 = A[25] & B[35];
    assign stage0_r26_c34 = A[26] & B[34];
    assign stage0_r27_c33 = A[27] & B[33];
    assign stage0_r28_c32 = A[28] & B[32];
    assign stage0_r29_c31 = A[29] & B[31];
    assign stage0_r30_c30 = A[30] & B[30];
    assign stage0_r31_c29 = A[31] & B[29];
    assign stage0_r32_c28 = A[32] & B[28];
    assign stage0_r33_c27 = A[33] & B[27];
    assign stage0_r34_c26 = A[34] & B[26];
    assign stage0_r35_c25 = A[35] & B[25];
    assign stage0_r36_c24 = A[36] & B[24];
    assign stage0_r37_c23 = A[37] & B[23];
    assign stage0_r38_c22 = A[38] & B[22];
    assign stage0_r39_c21 = A[39] & B[21];
    assign stage0_r40_c20 = A[40] & B[20];
    assign stage0_r41_c19 = A[41] & B[19];
    assign stage0_r42_c18 = A[42] & B[18];
    assign stage0_r43_c17 = A[43] & B[17];
    assign stage0_r44_c16 = A[44] & B[16];
    assign stage0_r45_c15 = A[45] & B[15];
    assign stage0_r46_c14 = A[46] & B[14];
    assign stage0_r47_c13 = A[47] & B[13];
    assign stage0_r48_c12 = A[48] & B[12];
    assign stage0_r49_c11 = A[49] & B[11];
    assign stage0_r50_c10 = A[50] & B[10];
    assign stage0_r51_c9 = A[51] & B[9];
    assign stage0_r52_c8 = A[52] & B[8];
    assign stage0_r53_c7 = A[53] & B[7];
    assign stage0_r54_c6 = A[54] & B[6];
    assign stage0_r55_c5 = A[55] & B[5];
    assign stage0_r56_c4 = A[56] & B[4];
    assign stage0_r57_c3 = A[57] & B[3];
    assign stage0_r58_c2 = A[58] & B[2];
    assign stage0_r59_c1 = A[59] & B[1];
    assign stage0_r60_c0 = A[60] & B[0];
    assign stage0_r21_c40 = A[21] & B[40];
    assign stage0_r22_c39 = A[22] & B[39];
    assign stage0_r23_c38 = A[23] & B[38];
    assign stage0_r24_c37 = A[24] & B[37];
    assign stage0_r25_c36 = A[25] & B[36];
    assign stage0_r26_c35 = A[26] & B[35];
    assign stage0_r27_c34 = A[27] & B[34];
    assign stage0_r28_c33 = A[28] & B[33];
    assign stage0_r29_c32 = A[29] & B[32];
    assign stage0_r30_c31 = A[30] & B[31];
    assign stage0_r31_c30 = A[31] & B[30];
    assign stage0_r32_c29 = A[32] & B[29];
    assign stage0_r33_c28 = A[33] & B[28];
    assign stage0_r34_c27 = A[34] & B[27];
    assign stage0_r35_c26 = A[35] & B[26];
    assign stage0_r36_c25 = A[36] & B[25];
    assign stage0_r37_c24 = A[37] & B[24];
    assign stage0_r38_c23 = A[38] & B[23];
    assign stage0_r39_c22 = A[39] & B[22];
    assign stage0_r40_c21 = A[40] & B[21];
    assign stage0_r41_c20 = A[41] & B[20];
    assign stage0_r42_c19 = A[42] & B[19];
    assign stage0_r43_c18 = A[43] & B[18];
    assign stage0_r44_c17 = A[44] & B[17];
    assign stage0_r45_c16 = A[45] & B[16];
    assign stage0_r46_c15 = A[46] & B[15];
    assign stage0_r47_c14 = A[47] & B[14];
    assign stage0_r48_c13 = A[48] & B[13];
    assign stage0_r49_c12 = A[49] & B[12];
    assign stage0_r50_c11 = A[50] & B[11];
    assign stage0_r51_c10 = A[51] & B[10];
    assign stage0_r52_c9 = A[52] & B[9];
    assign stage0_r53_c8 = A[53] & B[8];
    assign stage0_r54_c7 = A[54] & B[7];
    assign stage0_r55_c6 = A[55] & B[6];
    assign stage0_r56_c5 = A[56] & B[5];
    assign stage0_r57_c4 = A[57] & B[4];
    assign stage0_r58_c3 = A[58] & B[3];
    assign stage0_r59_c2 = A[59] & B[2];
    assign stage0_r60_c1 = A[60] & B[1];
    assign stage0_r61_c0 = A[61] & B[0];
    assign stage0_r22_c40 = A[22] & B[40];
    assign stage0_r23_c39 = A[23] & B[39];
    assign stage0_r24_c38 = A[24] & B[38];
    assign stage0_r25_c37 = A[25] & B[37];
    assign stage0_r26_c36 = A[26] & B[36];
    assign stage0_r27_c35 = A[27] & B[35];
    assign stage0_r28_c34 = A[28] & B[34];
    assign stage0_r29_c33 = A[29] & B[33];
    assign stage0_r30_c32 = A[30] & B[32];
    assign stage0_r31_c31 = A[31] & B[31];
    assign stage0_r32_c30 = A[32] & B[30];
    assign stage0_r33_c29 = A[33] & B[29];
    assign stage0_r34_c28 = A[34] & B[28];
    assign stage0_r35_c27 = A[35] & B[27];
    assign stage0_r36_c26 = A[36] & B[26];
    assign stage0_r37_c25 = A[37] & B[25];
    assign stage0_r38_c24 = A[38] & B[24];
    assign stage0_r39_c23 = A[39] & B[23];
    assign stage0_r40_c22 = A[40] & B[22];
    assign stage0_r41_c21 = A[41] & B[21];
    assign stage0_r42_c20 = A[42] & B[20];
    assign stage0_r43_c19 = A[43] & B[19];
    assign stage0_r44_c18 = A[44] & B[18];
    assign stage0_r45_c17 = A[45] & B[17];
    assign stage0_r46_c16 = A[46] & B[16];
    assign stage0_r47_c15 = A[47] & B[15];
    assign stage0_r48_c14 = A[48] & B[14];
    assign stage0_r49_c13 = A[49] & B[13];
    assign stage0_r50_c12 = A[50] & B[12];
    assign stage0_r51_c11 = A[51] & B[11];
    assign stage0_r52_c10 = A[52] & B[10];
    assign stage0_r53_c9 = A[53] & B[9];
    assign stage0_r54_c8 = A[54] & B[8];
    assign stage0_r55_c7 = A[55] & B[7];
    assign stage0_r56_c6 = A[56] & B[6];
    assign stage0_r57_c5 = A[57] & B[5];
    assign stage0_r58_c4 = A[58] & B[4];
    assign stage0_r59_c3 = A[59] & B[3];
    assign stage0_r60_c2 = A[60] & B[2];
    assign stage0_r61_c1 = A[61] & B[1];
    assign stage0_r62_c0 = A[62] & B[0];
    assign stage0_r23_c40 = A[23] & B[40];
    assign stage0_r24_c39 = A[24] & B[39];
    assign stage0_r25_c38 = A[25] & B[38];
    assign stage0_r26_c37 = A[26] & B[37];
    assign stage0_r27_c36 = A[27] & B[36];
    assign stage0_r28_c35 = A[28] & B[35];
    assign stage0_r29_c34 = A[29] & B[34];
    assign stage0_r30_c33 = A[30] & B[33];
    assign stage0_r31_c32 = A[31] & B[32];
    assign stage0_r32_c31 = A[32] & B[31];
    assign stage0_r33_c30 = A[33] & B[30];
    assign stage0_r34_c29 = A[34] & B[29];
    assign stage0_r35_c28 = A[35] & B[28];
    assign stage0_r36_c27 = A[36] & B[27];
    assign stage0_r37_c26 = A[37] & B[26];
    assign stage0_r38_c25 = A[38] & B[25];
    assign stage0_r39_c24 = A[39] & B[24];
    assign stage0_r40_c23 = A[40] & B[23];
    assign stage0_r41_c22 = A[41] & B[22];
    assign stage0_r42_c21 = A[42] & B[21];
    assign stage0_r43_c20 = A[43] & B[20];
    assign stage0_r44_c19 = A[44] & B[19];
    assign stage0_r45_c18 = A[45] & B[18];
    assign stage0_r46_c17 = A[46] & B[17];
    assign stage0_r47_c16 = A[47] & B[16];
    assign stage0_r48_c15 = A[48] & B[15];
    assign stage0_r49_c14 = A[49] & B[14];
    assign stage0_r50_c13 = A[50] & B[13];
    assign stage0_r51_c12 = A[51] & B[12];
    assign stage0_r52_c11 = A[52] & B[11];
    assign stage0_r53_c10 = A[53] & B[10];
    assign stage0_r54_c9 = A[54] & B[9];
    assign stage0_r55_c8 = A[55] & B[8];
    assign stage0_r56_c7 = A[56] & B[7];
    assign stage0_r57_c6 = A[57] & B[6];
    assign stage0_r58_c5 = A[58] & B[5];
    assign stage0_r59_c4 = A[59] & B[4];
    assign stage0_r60_c3 = A[60] & B[3];
    assign stage0_r61_c2 = A[61] & B[2];
    assign stage0_r62_c1 = A[62] & B[1];
    assign stage0_r63_c0 = A[63] & B[0];
    assign stage0_r24_c40 = A[24] & B[40];
    assign stage0_r25_c39 = A[25] & B[39];
    assign stage0_r26_c38 = A[26] & B[38];
    assign stage0_r27_c37 = A[27] & B[37];
    assign stage0_r28_c36 = A[28] & B[36];
    assign stage0_r29_c35 = A[29] & B[35];
    assign stage0_r30_c34 = A[30] & B[34];
    assign stage0_r31_c33 = A[31] & B[33];
    assign stage0_r32_c32 = A[32] & B[32];
    assign stage0_r33_c31 = A[33] & B[31];
    assign stage0_r34_c30 = A[34] & B[30];
    assign stage0_r35_c29 = A[35] & B[29];
    assign stage0_r36_c28 = A[36] & B[28];
    assign stage0_r37_c27 = A[37] & B[27];
    assign stage0_r38_c26 = A[38] & B[26];
    assign stage0_r39_c25 = A[39] & B[25];
    assign stage0_r40_c24 = A[40] & B[24];
    assign stage0_r41_c23 = A[41] & B[23];
    assign stage0_r42_c22 = A[42] & B[22];
    assign stage0_r43_c21 = A[43] & B[21];
    assign stage0_r44_c20 = A[44] & B[20];
    assign stage0_r45_c19 = A[45] & B[19];
    assign stage0_r46_c18 = A[46] & B[18];
    assign stage0_r47_c17 = A[47] & B[17];
    assign stage0_r48_c16 = A[48] & B[16];
    assign stage0_r49_c15 = A[49] & B[15];
    assign stage0_r50_c14 = A[50] & B[14];
    assign stage0_r51_c13 = A[51] & B[13];
    assign stage0_r52_c12 = A[52] & B[12];
    assign stage0_r53_c11 = A[53] & B[11];
    assign stage0_r54_c10 = A[54] & B[10];
    assign stage0_r55_c9 = A[55] & B[9];
    assign stage0_r56_c8 = A[56] & B[8];
    assign stage0_r57_c7 = A[57] & B[7];
    assign stage0_r58_c6 = A[58] & B[6];
    assign stage0_r59_c5 = A[59] & B[5];
    assign stage0_r60_c4 = A[60] & B[4];
    assign stage0_r61_c3 = A[61] & B[3];
    assign stage0_r62_c2 = A[62] & B[2];
    assign stage0_r63_c1 = A[63] & B[1];
    assign stage0_r64_c0 = A[64] & B[0];
    assign stage0_r25_c40 = A[25] & B[40];
    assign stage0_r26_c39 = A[26] & B[39];
    assign stage0_r27_c38 = A[27] & B[38];
    assign stage0_r28_c37 = A[28] & B[37];
    assign stage0_r29_c36 = A[29] & B[36];
    assign stage0_r30_c35 = A[30] & B[35];
    assign stage0_r31_c34 = A[31] & B[34];
    assign stage0_r32_c33 = A[32] & B[33];
    assign stage0_r33_c32 = A[33] & B[32];
    assign stage0_r34_c31 = A[34] & B[31];
    assign stage0_r35_c30 = A[35] & B[30];
    assign stage0_r36_c29 = A[36] & B[29];
    assign stage0_r37_c28 = A[37] & B[28];
    assign stage0_r38_c27 = A[38] & B[27];
    assign stage0_r39_c26 = A[39] & B[26];
    assign stage0_r40_c25 = A[40] & B[25];
    assign stage0_r41_c24 = A[41] & B[24];
    assign stage0_r42_c23 = A[42] & B[23];
    assign stage0_r43_c22 = A[43] & B[22];
    assign stage0_r44_c21 = A[44] & B[21];
    assign stage0_r45_c20 = A[45] & B[20];
    assign stage0_r46_c19 = A[46] & B[19];
    assign stage0_r47_c18 = A[47] & B[18];
    assign stage0_r48_c17 = A[48] & B[17];
    assign stage0_r49_c16 = A[49] & B[16];
    assign stage0_r50_c15 = A[50] & B[15];
    assign stage0_r51_c14 = A[51] & B[14];
    assign stage0_r52_c13 = A[52] & B[13];
    assign stage0_r53_c12 = A[53] & B[12];
    assign stage0_r54_c11 = A[54] & B[11];
    assign stage0_r55_c10 = A[55] & B[10];
    assign stage0_r56_c9 = A[56] & B[9];
    assign stage0_r57_c8 = A[57] & B[8];
    assign stage0_r58_c7 = A[58] & B[7];
    assign stage0_r59_c6 = A[59] & B[6];
    assign stage0_r60_c5 = A[60] & B[5];
    assign stage0_r61_c4 = A[61] & B[4];
    assign stage0_r62_c3 = A[62] & B[3];
    assign stage0_r63_c2 = A[63] & B[2];
    assign stage0_r64_c1 = A[64] & B[1];
    assign stage0_r65_c0 = A[65] & B[0];
    assign stage0_r26_c40 = A[26] & B[40];
    assign stage0_r27_c39 = A[27] & B[39];
    assign stage0_r28_c38 = A[28] & B[38];
    assign stage0_r29_c37 = A[29] & B[37];
    assign stage0_r30_c36 = A[30] & B[36];
    assign stage0_r31_c35 = A[31] & B[35];
    assign stage0_r32_c34 = A[32] & B[34];
    assign stage0_r33_c33 = A[33] & B[33];
    assign stage0_r34_c32 = A[34] & B[32];
    assign stage0_r35_c31 = A[35] & B[31];
    assign stage0_r36_c30 = A[36] & B[30];
    assign stage0_r37_c29 = A[37] & B[29];
    assign stage0_r38_c28 = A[38] & B[28];
    assign stage0_r39_c27 = A[39] & B[27];
    assign stage0_r40_c26 = A[40] & B[26];
    assign stage0_r41_c25 = A[41] & B[25];
    assign stage0_r42_c24 = A[42] & B[24];
    assign stage0_r43_c23 = A[43] & B[23];
    assign stage0_r44_c22 = A[44] & B[22];
    assign stage0_r45_c21 = A[45] & B[21];
    assign stage0_r46_c20 = A[46] & B[20];
    assign stage0_r47_c19 = A[47] & B[19];
    assign stage0_r48_c18 = A[48] & B[18];
    assign stage0_r49_c17 = A[49] & B[17];
    assign stage0_r50_c16 = A[50] & B[16];
    assign stage0_r51_c15 = A[51] & B[15];
    assign stage0_r52_c14 = A[52] & B[14];
    assign stage0_r53_c13 = A[53] & B[13];
    assign stage0_r54_c12 = A[54] & B[12];
    assign stage0_r55_c11 = A[55] & B[11];
    assign stage0_r56_c10 = A[56] & B[10];
    assign stage0_r57_c9 = A[57] & B[9];
    assign stage0_r58_c8 = A[58] & B[8];
    assign stage0_r59_c7 = A[59] & B[7];
    assign stage0_r60_c6 = A[60] & B[6];
    assign stage0_r61_c5 = A[61] & B[5];
    assign stage0_r62_c4 = A[62] & B[4];
    assign stage0_r63_c3 = A[63] & B[3];
    assign stage0_r64_c2 = A[64] & B[2];
    assign stage0_r65_c1 = A[65] & B[1];
    assign stage0_r66_c0 = A[66] & B[0];
    assign stage0_r27_c40 = A[27] & B[40];
    assign stage0_r28_c39 = A[28] & B[39];
    assign stage0_r29_c38 = A[29] & B[38];
    assign stage0_r30_c37 = A[30] & B[37];
    assign stage0_r31_c36 = A[31] & B[36];
    assign stage0_r32_c35 = A[32] & B[35];
    assign stage0_r33_c34 = A[33] & B[34];
    assign stage0_r34_c33 = A[34] & B[33];
    assign stage0_r35_c32 = A[35] & B[32];
    assign stage0_r36_c31 = A[36] & B[31];
    assign stage0_r37_c30 = A[37] & B[30];
    assign stage0_r38_c29 = A[38] & B[29];
    assign stage0_r39_c28 = A[39] & B[28];
    assign stage0_r40_c27 = A[40] & B[27];
    assign stage0_r41_c26 = A[41] & B[26];
    assign stage0_r42_c25 = A[42] & B[25];
    assign stage0_r43_c24 = A[43] & B[24];
    assign stage0_r44_c23 = A[44] & B[23];
    assign stage0_r45_c22 = A[45] & B[22];
    assign stage0_r46_c21 = A[46] & B[21];
    assign stage0_r47_c20 = A[47] & B[20];
    assign stage0_r48_c19 = A[48] & B[19];
    assign stage0_r49_c18 = A[49] & B[18];
    assign stage0_r50_c17 = A[50] & B[17];
    assign stage0_r51_c16 = A[51] & B[16];
    assign stage0_r52_c15 = A[52] & B[15];
    assign stage0_r53_c14 = A[53] & B[14];
    assign stage0_r54_c13 = A[54] & B[13];
    assign stage0_r55_c12 = A[55] & B[12];
    assign stage0_r56_c11 = A[56] & B[11];
    assign stage0_r57_c10 = A[57] & B[10];
    assign stage0_r58_c9 = A[58] & B[9];
    assign stage0_r59_c8 = A[59] & B[8];
    assign stage0_r60_c7 = A[60] & B[7];
    assign stage0_r61_c6 = A[61] & B[6];
    assign stage0_r62_c5 = A[62] & B[5];
    assign stage0_r63_c4 = A[63] & B[4];
    assign stage0_r64_c3 = A[64] & B[3];
    assign stage0_r65_c2 = A[65] & B[2];
    assign stage0_r66_c1 = A[66] & B[1];
    assign stage0_r67_c0 = A[67] & B[0];
    assign stage0_r28_c40 = A[28] & B[40];
    assign stage0_r29_c39 = A[29] & B[39];
    assign stage0_r30_c38 = A[30] & B[38];
    assign stage0_r31_c37 = A[31] & B[37];
    assign stage0_r32_c36 = A[32] & B[36];
    assign stage0_r33_c35 = A[33] & B[35];
    assign stage0_r34_c34 = A[34] & B[34];
    assign stage0_r35_c33 = A[35] & B[33];
    assign stage0_r36_c32 = A[36] & B[32];
    assign stage0_r37_c31 = A[37] & B[31];
    assign stage0_r38_c30 = A[38] & B[30];
    assign stage0_r39_c29 = A[39] & B[29];
    assign stage0_r40_c28 = A[40] & B[28];
    assign stage0_r41_c27 = A[41] & B[27];
    assign stage0_r42_c26 = A[42] & B[26];
    assign stage0_r43_c25 = A[43] & B[25];
    assign stage0_r44_c24 = A[44] & B[24];
    assign stage0_r45_c23 = A[45] & B[23];
    assign stage0_r46_c22 = A[46] & B[22];
    assign stage0_r47_c21 = A[47] & B[21];
    assign stage0_r48_c20 = A[48] & B[20];
    assign stage0_r49_c19 = A[49] & B[19];
    assign stage0_r50_c18 = A[50] & B[18];
    assign stage0_r51_c17 = A[51] & B[17];
    assign stage0_r52_c16 = A[52] & B[16];
    assign stage0_r53_c15 = A[53] & B[15];
    assign stage0_r54_c14 = A[54] & B[14];
    assign stage0_r55_c13 = A[55] & B[13];
    assign stage0_r56_c12 = A[56] & B[12];
    assign stage0_r57_c11 = A[57] & B[11];
    assign stage0_r58_c10 = A[58] & B[10];
    assign stage0_r59_c9 = A[59] & B[9];
    assign stage0_r60_c8 = A[60] & B[8];
    assign stage0_r61_c7 = A[61] & B[7];
    assign stage0_r62_c6 = A[62] & B[6];
    assign stage0_r63_c5 = A[63] & B[5];
    assign stage0_r64_c4 = A[64] & B[4];
    assign stage0_r65_c3 = A[65] & B[3];
    assign stage0_r66_c2 = A[66] & B[2];
    assign stage0_r67_c1 = A[67] & B[1];
    assign stage0_r68_c0 = A[68] & B[0];
    assign stage0_r29_c40 = A[29] & B[40];
    assign stage0_r30_c39 = A[30] & B[39];
    assign stage0_r31_c38 = A[31] & B[38];
    assign stage0_r32_c37 = A[32] & B[37];
    assign stage0_r33_c36 = A[33] & B[36];
    assign stage0_r34_c35 = A[34] & B[35];
    assign stage0_r35_c34 = A[35] & B[34];
    assign stage0_r36_c33 = A[36] & B[33];
    assign stage0_r37_c32 = A[37] & B[32];
    assign stage0_r38_c31 = A[38] & B[31];
    assign stage0_r39_c30 = A[39] & B[30];
    assign stage0_r40_c29 = A[40] & B[29];
    assign stage0_r41_c28 = A[41] & B[28];
    assign stage0_r42_c27 = A[42] & B[27];
    assign stage0_r43_c26 = A[43] & B[26];
    assign stage0_r44_c25 = A[44] & B[25];
    assign stage0_r45_c24 = A[45] & B[24];
    assign stage0_r46_c23 = A[46] & B[23];
    assign stage0_r47_c22 = A[47] & B[22];
    assign stage0_r48_c21 = A[48] & B[21];
    assign stage0_r49_c20 = A[49] & B[20];
    assign stage0_r50_c19 = A[50] & B[19];
    assign stage0_r51_c18 = A[51] & B[18];
    assign stage0_r52_c17 = A[52] & B[17];
    assign stage0_r53_c16 = A[53] & B[16];
    assign stage0_r54_c15 = A[54] & B[15];
    assign stage0_r55_c14 = A[55] & B[14];
    assign stage0_r56_c13 = A[56] & B[13];
    assign stage0_r57_c12 = A[57] & B[12];
    assign stage0_r58_c11 = A[58] & B[11];
    assign stage0_r59_c10 = A[59] & B[10];
    assign stage0_r60_c9 = A[60] & B[9];
    assign stage0_r61_c8 = A[61] & B[8];
    assign stage0_r62_c7 = A[62] & B[7];
    assign stage0_r63_c6 = A[63] & B[6];
    assign stage0_r64_c5 = A[64] & B[5];
    assign stage0_r65_c4 = A[65] & B[4];
    assign stage0_r66_c3 = A[66] & B[3];
    assign stage0_r67_c2 = A[67] & B[2];
    assign stage0_r68_c1 = A[68] & B[1];
    assign stage0_r69_c0 = A[69] & B[0];
    assign stage0_r30_c40 = A[30] & B[40];
    assign stage0_r31_c39 = A[31] & B[39];
    assign stage0_r32_c38 = A[32] & B[38];
    assign stage0_r33_c37 = A[33] & B[37];
    assign stage0_r34_c36 = A[34] & B[36];
    assign stage0_r35_c35 = A[35] & B[35];
    assign stage0_r36_c34 = A[36] & B[34];
    assign stage0_r37_c33 = A[37] & B[33];
    assign stage0_r38_c32 = A[38] & B[32];
    assign stage0_r39_c31 = A[39] & B[31];
    assign stage0_r40_c30 = A[40] & B[30];
    assign stage0_r41_c29 = A[41] & B[29];
    assign stage0_r42_c28 = A[42] & B[28];
    assign stage0_r43_c27 = A[43] & B[27];
    assign stage0_r44_c26 = A[44] & B[26];
    assign stage0_r45_c25 = A[45] & B[25];
    assign stage0_r46_c24 = A[46] & B[24];
    assign stage0_r47_c23 = A[47] & B[23];
    assign stage0_r48_c22 = A[48] & B[22];
    assign stage0_r49_c21 = A[49] & B[21];
    assign stage0_r50_c20 = A[50] & B[20];
    assign stage0_r51_c19 = A[51] & B[19];
    assign stage0_r52_c18 = A[52] & B[18];
    assign stage0_r53_c17 = A[53] & B[17];
    assign stage0_r54_c16 = A[54] & B[16];
    assign stage0_r55_c15 = A[55] & B[15];
    assign stage0_r56_c14 = A[56] & B[14];
    assign stage0_r57_c13 = A[57] & B[13];
    assign stage0_r58_c12 = A[58] & B[12];
    assign stage0_r59_c11 = A[59] & B[11];
    assign stage0_r60_c10 = A[60] & B[10];
    assign stage0_r61_c9 = A[61] & B[9];
    assign stage0_r62_c8 = A[62] & B[8];
    assign stage0_r63_c7 = A[63] & B[7];
    assign stage0_r64_c6 = A[64] & B[6];
    assign stage0_r65_c5 = A[65] & B[5];
    assign stage0_r66_c4 = A[66] & B[4];
    assign stage0_r67_c3 = A[67] & B[3];
    assign stage0_r68_c2 = A[68] & B[2];
    assign stage0_r69_c1 = A[69] & B[1];
    assign stage0_r70_c0 = A[70] & B[0];
    assign stage0_r31_c40 = A[31] & B[40];
    assign stage0_r32_c39 = A[32] & B[39];
    assign stage0_r33_c38 = A[33] & B[38];
    assign stage0_r34_c37 = A[34] & B[37];
    assign stage0_r35_c36 = A[35] & B[36];
    assign stage0_r36_c35 = A[36] & B[35];
    assign stage0_r37_c34 = A[37] & B[34];
    assign stage0_r38_c33 = A[38] & B[33];
    assign stage0_r39_c32 = A[39] & B[32];
    assign stage0_r40_c31 = A[40] & B[31];
    assign stage0_r41_c30 = A[41] & B[30];
    assign stage0_r42_c29 = A[42] & B[29];
    assign stage0_r43_c28 = A[43] & B[28];
    assign stage0_r44_c27 = A[44] & B[27];
    assign stage0_r45_c26 = A[45] & B[26];
    assign stage0_r46_c25 = A[46] & B[25];
    assign stage0_r47_c24 = A[47] & B[24];
    assign stage0_r48_c23 = A[48] & B[23];
    assign stage0_r49_c22 = A[49] & B[22];
    assign stage0_r50_c21 = A[50] & B[21];
    assign stage0_r51_c20 = A[51] & B[20];
    assign stage0_r52_c19 = A[52] & B[19];
    assign stage0_r53_c18 = A[53] & B[18];
    assign stage0_r54_c17 = A[54] & B[17];
    assign stage0_r55_c16 = A[55] & B[16];
    assign stage0_r56_c15 = A[56] & B[15];
    assign stage0_r57_c14 = A[57] & B[14];
    assign stage0_r58_c13 = A[58] & B[13];
    assign stage0_r59_c12 = A[59] & B[12];
    assign stage0_r60_c11 = A[60] & B[11];
    assign stage0_r61_c10 = A[61] & B[10];
    assign stage0_r62_c9 = A[62] & B[9];
    assign stage0_r63_c8 = A[63] & B[8];
    assign stage0_r64_c7 = A[64] & B[7];
    assign stage0_r65_c6 = A[65] & B[6];
    assign stage0_r66_c5 = A[66] & B[5];
    assign stage0_r67_c4 = A[67] & B[4];
    assign stage0_r68_c3 = A[68] & B[3];
    assign stage0_r69_c2 = A[69] & B[2];
    assign stage0_r70_c1 = A[70] & B[1];
    assign stage0_r71_c0 = A[71] & B[0];
    assign stage0_r32_c40 = A[32] & B[40];
    assign stage0_r33_c39 = A[33] & B[39];
    assign stage0_r34_c38 = A[34] & B[38];
    assign stage0_r35_c37 = A[35] & B[37];
    assign stage0_r36_c36 = A[36] & B[36];
    assign stage0_r37_c35 = A[37] & B[35];
    assign stage0_r38_c34 = A[38] & B[34];
    assign stage0_r39_c33 = A[39] & B[33];
    assign stage0_r40_c32 = A[40] & B[32];
    assign stage0_r41_c31 = A[41] & B[31];
    assign stage0_r42_c30 = A[42] & B[30];
    assign stage0_r43_c29 = A[43] & B[29];
    assign stage0_r44_c28 = A[44] & B[28];
    assign stage0_r45_c27 = A[45] & B[27];
    assign stage0_r46_c26 = A[46] & B[26];
    assign stage0_r47_c25 = A[47] & B[25];
    assign stage0_r48_c24 = A[48] & B[24];
    assign stage0_r49_c23 = A[49] & B[23];
    assign stage0_r50_c22 = A[50] & B[22];
    assign stage0_r51_c21 = A[51] & B[21];
    assign stage0_r52_c20 = A[52] & B[20];
    assign stage0_r53_c19 = A[53] & B[19];
    assign stage0_r54_c18 = A[54] & B[18];
    assign stage0_r55_c17 = A[55] & B[17];
    assign stage0_r56_c16 = A[56] & B[16];
    assign stage0_r57_c15 = A[57] & B[15];
    assign stage0_r58_c14 = A[58] & B[14];
    assign stage0_r59_c13 = A[59] & B[13];
    assign stage0_r60_c12 = A[60] & B[12];
    assign stage0_r61_c11 = A[61] & B[11];
    assign stage0_r62_c10 = A[62] & B[10];
    assign stage0_r63_c9 = A[63] & B[9];
    assign stage0_r64_c8 = A[64] & B[8];
    assign stage0_r65_c7 = A[65] & B[7];
    assign stage0_r66_c6 = A[66] & B[6];
    assign stage0_r67_c5 = A[67] & B[5];
    assign stage0_r68_c4 = A[68] & B[4];
    assign stage0_r69_c3 = A[69] & B[3];
    assign stage0_r70_c2 = A[70] & B[2];
    assign stage0_r71_c1 = A[71] & B[1];
    assign stage0_r33_c40 = A[33] & B[40];
    assign stage0_r34_c39 = A[34] & B[39];
    assign stage0_r35_c38 = A[35] & B[38];
    assign stage0_r36_c37 = A[36] & B[37];
    assign stage0_r37_c36 = A[37] & B[36];
    assign stage0_r38_c35 = A[38] & B[35];
    assign stage0_r39_c34 = A[39] & B[34];
    assign stage0_r40_c33 = A[40] & B[33];
    assign stage0_r41_c32 = A[41] & B[32];
    assign stage0_r42_c31 = A[42] & B[31];
    assign stage0_r43_c30 = A[43] & B[30];
    assign stage0_r44_c29 = A[44] & B[29];
    assign stage0_r45_c28 = A[45] & B[28];
    assign stage0_r46_c27 = A[46] & B[27];
    assign stage0_r47_c26 = A[47] & B[26];
    assign stage0_r48_c25 = A[48] & B[25];
    assign stage0_r49_c24 = A[49] & B[24];
    assign stage0_r50_c23 = A[50] & B[23];
    assign stage0_r51_c22 = A[51] & B[22];
    assign stage0_r52_c21 = A[52] & B[21];
    assign stage0_r53_c20 = A[53] & B[20];
    assign stage0_r54_c19 = A[54] & B[19];
    assign stage0_r55_c18 = A[55] & B[18];
    assign stage0_r56_c17 = A[56] & B[17];
    assign stage0_r57_c16 = A[57] & B[16];
    assign stage0_r58_c15 = A[58] & B[15];
    assign stage0_r59_c14 = A[59] & B[14];
    assign stage0_r60_c13 = A[60] & B[13];
    assign stage0_r61_c12 = A[61] & B[12];
    assign stage0_r62_c11 = A[62] & B[11];
    assign stage0_r63_c10 = A[63] & B[10];
    assign stage0_r64_c9 = A[64] & B[9];
    assign stage0_r65_c8 = A[65] & B[8];
    assign stage0_r66_c7 = A[66] & B[7];
    assign stage0_r67_c6 = A[67] & B[6];
    assign stage0_r68_c5 = A[68] & B[5];
    assign stage0_r69_c4 = A[69] & B[4];
    assign stage0_r70_c3 = A[70] & B[3];
    assign stage0_r71_c2 = A[71] & B[2];
    assign stage0_r34_c40 = A[34] & B[40];
    assign stage0_r35_c39 = A[35] & B[39];
    assign stage0_r36_c38 = A[36] & B[38];
    assign stage0_r37_c37 = A[37] & B[37];
    assign stage0_r38_c36 = A[38] & B[36];
    assign stage0_r39_c35 = A[39] & B[35];
    assign stage0_r40_c34 = A[40] & B[34];
    assign stage0_r41_c33 = A[41] & B[33];
    assign stage0_r42_c32 = A[42] & B[32];
    assign stage0_r43_c31 = A[43] & B[31];
    assign stage0_r44_c30 = A[44] & B[30];
    assign stage0_r45_c29 = A[45] & B[29];
    assign stage0_r46_c28 = A[46] & B[28];
    assign stage0_r47_c27 = A[47] & B[27];
    assign stage0_r48_c26 = A[48] & B[26];
    assign stage0_r49_c25 = A[49] & B[25];
    assign stage0_r50_c24 = A[50] & B[24];
    assign stage0_r51_c23 = A[51] & B[23];
    assign stage0_r52_c22 = A[52] & B[22];
    assign stage0_r53_c21 = A[53] & B[21];
    assign stage0_r54_c20 = A[54] & B[20];
    assign stage0_r55_c19 = A[55] & B[19];
    assign stage0_r56_c18 = A[56] & B[18];
    assign stage0_r57_c17 = A[57] & B[17];
    assign stage0_r58_c16 = A[58] & B[16];
    assign stage0_r59_c15 = A[59] & B[15];
    assign stage0_r60_c14 = A[60] & B[14];
    assign stage0_r61_c13 = A[61] & B[13];
    assign stage0_r62_c12 = A[62] & B[12];
    assign stage0_r63_c11 = A[63] & B[11];
    assign stage0_r64_c10 = A[64] & B[10];
    assign stage0_r65_c9 = A[65] & B[9];
    assign stage0_r66_c8 = A[66] & B[8];
    assign stage0_r67_c7 = A[67] & B[7];
    assign stage0_r68_c6 = A[68] & B[6];
    assign stage0_r69_c5 = A[69] & B[5];
    assign stage0_r70_c4 = A[70] & B[4];
    assign stage0_r71_c3 = A[71] & B[3];
    assign stage0_r35_c40 = A[35] & B[40];
    assign stage0_r36_c39 = A[36] & B[39];
    assign stage0_r37_c38 = A[37] & B[38];
    assign stage0_r38_c37 = A[38] & B[37];
    assign stage0_r39_c36 = A[39] & B[36];
    assign stage0_r40_c35 = A[40] & B[35];
    assign stage0_r41_c34 = A[41] & B[34];
    assign stage0_r42_c33 = A[42] & B[33];
    assign stage0_r43_c32 = A[43] & B[32];
    assign stage0_r44_c31 = A[44] & B[31];
    assign stage0_r45_c30 = A[45] & B[30];
    assign stage0_r46_c29 = A[46] & B[29];
    assign stage0_r47_c28 = A[47] & B[28];
    assign stage0_r48_c27 = A[48] & B[27];
    assign stage0_r49_c26 = A[49] & B[26];
    assign stage0_r50_c25 = A[50] & B[25];
    assign stage0_r51_c24 = A[51] & B[24];
    assign stage0_r52_c23 = A[52] & B[23];
    assign stage0_r53_c22 = A[53] & B[22];
    assign stage0_r54_c21 = A[54] & B[21];
    assign stage0_r55_c20 = A[55] & B[20];
    assign stage0_r56_c19 = A[56] & B[19];
    assign stage0_r57_c18 = A[57] & B[18];
    assign stage0_r58_c17 = A[58] & B[17];
    assign stage0_r59_c16 = A[59] & B[16];
    assign stage0_r60_c15 = A[60] & B[15];
    assign stage0_r61_c14 = A[61] & B[14];
    assign stage0_r62_c13 = A[62] & B[13];
    assign stage0_r63_c12 = A[63] & B[12];
    assign stage0_r64_c11 = A[64] & B[11];
    assign stage0_r65_c10 = A[65] & B[10];
    assign stage0_r66_c9 = A[66] & B[9];
    assign stage0_r67_c8 = A[67] & B[8];
    assign stage0_r68_c7 = A[68] & B[7];
    assign stage0_r69_c6 = A[69] & B[6];
    assign stage0_r70_c5 = A[70] & B[5];
    assign stage0_r71_c4 = A[71] & B[4];
    assign stage0_r36_c40 = A[36] & B[40];
    assign stage0_r37_c39 = A[37] & B[39];
    assign stage0_r38_c38 = A[38] & B[38];
    assign stage0_r39_c37 = A[39] & B[37];
    assign stage0_r40_c36 = A[40] & B[36];
    assign stage0_r41_c35 = A[41] & B[35];
    assign stage0_r42_c34 = A[42] & B[34];
    assign stage0_r43_c33 = A[43] & B[33];
    assign stage0_r44_c32 = A[44] & B[32];
    assign stage0_r45_c31 = A[45] & B[31];
    assign stage0_r46_c30 = A[46] & B[30];
    assign stage0_r47_c29 = A[47] & B[29];
    assign stage0_r48_c28 = A[48] & B[28];
    assign stage0_r49_c27 = A[49] & B[27];
    assign stage0_r50_c26 = A[50] & B[26];
    assign stage0_r51_c25 = A[51] & B[25];
    assign stage0_r52_c24 = A[52] & B[24];
    assign stage0_r53_c23 = A[53] & B[23];
    assign stage0_r54_c22 = A[54] & B[22];
    assign stage0_r55_c21 = A[55] & B[21];
    assign stage0_r56_c20 = A[56] & B[20];
    assign stage0_r57_c19 = A[57] & B[19];
    assign stage0_r58_c18 = A[58] & B[18];
    assign stage0_r59_c17 = A[59] & B[17];
    assign stage0_r60_c16 = A[60] & B[16];
    assign stage0_r61_c15 = A[61] & B[15];
    assign stage0_r62_c14 = A[62] & B[14];
    assign stage0_r63_c13 = A[63] & B[13];
    assign stage0_r64_c12 = A[64] & B[12];
    assign stage0_r65_c11 = A[65] & B[11];
    assign stage0_r66_c10 = A[66] & B[10];
    assign stage0_r67_c9 = A[67] & B[9];
    assign stage0_r68_c8 = A[68] & B[8];
    assign stage0_r69_c7 = A[69] & B[7];
    assign stage0_r70_c6 = A[70] & B[6];
    assign stage0_r71_c5 = A[71] & B[5];
    assign stage0_r37_c40 = A[37] & B[40];
    assign stage0_r38_c39 = A[38] & B[39];
    assign stage0_r39_c38 = A[39] & B[38];
    assign stage0_r40_c37 = A[40] & B[37];
    assign stage0_r41_c36 = A[41] & B[36];
    assign stage0_r42_c35 = A[42] & B[35];
    assign stage0_r43_c34 = A[43] & B[34];
    assign stage0_r44_c33 = A[44] & B[33];
    assign stage0_r45_c32 = A[45] & B[32];
    assign stage0_r46_c31 = A[46] & B[31];
    assign stage0_r47_c30 = A[47] & B[30];
    assign stage0_r48_c29 = A[48] & B[29];
    assign stage0_r49_c28 = A[49] & B[28];
    assign stage0_r50_c27 = A[50] & B[27];
    assign stage0_r51_c26 = A[51] & B[26];
    assign stage0_r52_c25 = A[52] & B[25];
    assign stage0_r53_c24 = A[53] & B[24];
    assign stage0_r54_c23 = A[54] & B[23];
    assign stage0_r55_c22 = A[55] & B[22];
    assign stage0_r56_c21 = A[56] & B[21];
    assign stage0_r57_c20 = A[57] & B[20];
    assign stage0_r58_c19 = A[58] & B[19];
    assign stage0_r59_c18 = A[59] & B[18];
    assign stage0_r60_c17 = A[60] & B[17];
    assign stage0_r61_c16 = A[61] & B[16];
    assign stage0_r62_c15 = A[62] & B[15];
    assign stage0_r63_c14 = A[63] & B[14];
    assign stage0_r64_c13 = A[64] & B[13];
    assign stage0_r65_c12 = A[65] & B[12];
    assign stage0_r66_c11 = A[66] & B[11];
    assign stage0_r67_c10 = A[67] & B[10];
    assign stage0_r68_c9 = A[68] & B[9];
    assign stage0_r69_c8 = A[69] & B[8];
    assign stage0_r70_c7 = A[70] & B[7];
    assign stage0_r71_c6 = A[71] & B[6];
    assign stage0_r38_c40 = A[38] & B[40];
    assign stage0_r39_c39 = A[39] & B[39];
    assign stage0_r40_c38 = A[40] & B[38];
    assign stage0_r41_c37 = A[41] & B[37];
    assign stage0_r42_c36 = A[42] & B[36];
    assign stage0_r43_c35 = A[43] & B[35];
    assign stage0_r44_c34 = A[44] & B[34];
    assign stage0_r45_c33 = A[45] & B[33];
    assign stage0_r46_c32 = A[46] & B[32];
    assign stage0_r47_c31 = A[47] & B[31];
    assign stage0_r48_c30 = A[48] & B[30];
    assign stage0_r49_c29 = A[49] & B[29];
    assign stage0_r50_c28 = A[50] & B[28];
    assign stage0_r51_c27 = A[51] & B[27];
    assign stage0_r52_c26 = A[52] & B[26];
    assign stage0_r53_c25 = A[53] & B[25];
    assign stage0_r54_c24 = A[54] & B[24];
    assign stage0_r55_c23 = A[55] & B[23];
    assign stage0_r56_c22 = A[56] & B[22];
    assign stage0_r57_c21 = A[57] & B[21];
    assign stage0_r58_c20 = A[58] & B[20];
    assign stage0_r59_c19 = A[59] & B[19];
    assign stage0_r60_c18 = A[60] & B[18];
    assign stage0_r61_c17 = A[61] & B[17];
    assign stage0_r62_c16 = A[62] & B[16];
    assign stage0_r63_c15 = A[63] & B[15];
    assign stage0_r64_c14 = A[64] & B[14];
    assign stage0_r65_c13 = A[65] & B[13];
    assign stage0_r66_c12 = A[66] & B[12];
    assign stage0_r67_c11 = A[67] & B[11];
    assign stage0_r68_c10 = A[68] & B[10];
    assign stage0_r69_c9 = A[69] & B[9];
    assign stage0_r70_c8 = A[70] & B[8];
    assign stage0_r71_c7 = A[71] & B[7];
    assign stage0_r39_c40 = A[39] & B[40];
    assign stage0_r40_c39 = A[40] & B[39];
    assign stage0_r41_c38 = A[41] & B[38];
    assign stage0_r42_c37 = A[42] & B[37];
    assign stage0_r43_c36 = A[43] & B[36];
    assign stage0_r44_c35 = A[44] & B[35];
    assign stage0_r45_c34 = A[45] & B[34];
    assign stage0_r46_c33 = A[46] & B[33];
    assign stage0_r47_c32 = A[47] & B[32];
    assign stage0_r48_c31 = A[48] & B[31];
    assign stage0_r49_c30 = A[49] & B[30];
    assign stage0_r50_c29 = A[50] & B[29];
    assign stage0_r51_c28 = A[51] & B[28];
    assign stage0_r52_c27 = A[52] & B[27];
    assign stage0_r53_c26 = A[53] & B[26];
    assign stage0_r54_c25 = A[54] & B[25];
    assign stage0_r55_c24 = A[55] & B[24];
    assign stage0_r56_c23 = A[56] & B[23];
    assign stage0_r57_c22 = A[57] & B[22];
    assign stage0_r58_c21 = A[58] & B[21];
    assign stage0_r59_c20 = A[59] & B[20];
    assign stage0_r60_c19 = A[60] & B[19];
    assign stage0_r61_c18 = A[61] & B[18];
    assign stage0_r62_c17 = A[62] & B[17];
    assign stage0_r63_c16 = A[63] & B[16];
    assign stage0_r64_c15 = A[64] & B[15];
    assign stage0_r65_c14 = A[65] & B[14];
    assign stage0_r66_c13 = A[66] & B[13];
    assign stage0_r67_c12 = A[67] & B[12];
    assign stage0_r68_c11 = A[68] & B[11];
    assign stage0_r69_c10 = A[69] & B[10];
    assign stage0_r70_c9 = A[70] & B[9];
    assign stage0_r71_c8 = A[71] & B[8];
    assign stage0_r40_c40 = A[40] & B[40];
    assign stage0_r41_c39 = A[41] & B[39];
    assign stage0_r42_c38 = A[42] & B[38];
    assign stage0_r43_c37 = A[43] & B[37];
    assign stage0_r44_c36 = A[44] & B[36];
    assign stage0_r45_c35 = A[45] & B[35];
    assign stage0_r46_c34 = A[46] & B[34];
    assign stage0_r47_c33 = A[47] & B[33];
    assign stage0_r48_c32 = A[48] & B[32];
    assign stage0_r49_c31 = A[49] & B[31];
    assign stage0_r50_c30 = A[50] & B[30];
    assign stage0_r51_c29 = A[51] & B[29];
    assign stage0_r52_c28 = A[52] & B[28];
    assign stage0_r53_c27 = A[53] & B[27];
    assign stage0_r54_c26 = A[54] & B[26];
    assign stage0_r55_c25 = A[55] & B[25];
    assign stage0_r56_c24 = A[56] & B[24];
    assign stage0_r57_c23 = A[57] & B[23];
    assign stage0_r58_c22 = A[58] & B[22];
    assign stage0_r59_c21 = A[59] & B[21];
    assign stage0_r60_c20 = A[60] & B[20];
    assign stage0_r61_c19 = A[61] & B[19];
    assign stage0_r62_c18 = A[62] & B[18];
    assign stage0_r63_c17 = A[63] & B[17];
    assign stage0_r64_c16 = A[64] & B[16];
    assign stage0_r65_c15 = A[65] & B[15];
    assign stage0_r66_c14 = A[66] & B[14];
    assign stage0_r67_c13 = A[67] & B[13];
    assign stage0_r68_c12 = A[68] & B[12];
    assign stage0_r69_c11 = A[69] & B[11];
    assign stage0_r70_c10 = A[70] & B[10];
    assign stage0_r71_c9 = A[71] & B[9];
    assign stage0_r41_c40 = A[41] & B[40];
    assign stage0_r42_c39 = A[42] & B[39];
    assign stage0_r43_c38 = A[43] & B[38];
    assign stage0_r44_c37 = A[44] & B[37];
    assign stage0_r45_c36 = A[45] & B[36];
    assign stage0_r46_c35 = A[46] & B[35];
    assign stage0_r47_c34 = A[47] & B[34];
    assign stage0_r48_c33 = A[48] & B[33];
    assign stage0_r49_c32 = A[49] & B[32];
    assign stage0_r50_c31 = A[50] & B[31];
    assign stage0_r51_c30 = A[51] & B[30];
    assign stage0_r52_c29 = A[52] & B[29];
    assign stage0_r53_c28 = A[53] & B[28];
    assign stage0_r54_c27 = A[54] & B[27];
    assign stage0_r55_c26 = A[55] & B[26];
    assign stage0_r56_c25 = A[56] & B[25];
    assign stage0_r57_c24 = A[57] & B[24];
    assign stage0_r58_c23 = A[58] & B[23];
    assign stage0_r59_c22 = A[59] & B[22];
    assign stage0_r60_c21 = A[60] & B[21];
    assign stage0_r61_c20 = A[61] & B[20];
    assign stage0_r62_c19 = A[62] & B[19];
    assign stage0_r63_c18 = A[63] & B[18];
    assign stage0_r64_c17 = A[64] & B[17];
    assign stage0_r65_c16 = A[65] & B[16];
    assign stage0_r66_c15 = A[66] & B[15];
    assign stage0_r67_c14 = A[67] & B[14];
    assign stage0_r68_c13 = A[68] & B[13];
    assign stage0_r69_c12 = A[69] & B[12];
    assign stage0_r70_c11 = A[70] & B[11];
    assign stage0_r71_c10 = A[71] & B[10];
    assign stage0_r42_c40 = A[42] & B[40];
    assign stage0_r43_c39 = A[43] & B[39];
    assign stage0_r44_c38 = A[44] & B[38];
    assign stage0_r45_c37 = A[45] & B[37];
    assign stage0_r46_c36 = A[46] & B[36];
    assign stage0_r47_c35 = A[47] & B[35];
    assign stage0_r48_c34 = A[48] & B[34];
    assign stage0_r49_c33 = A[49] & B[33];
    assign stage0_r50_c32 = A[50] & B[32];
    assign stage0_r51_c31 = A[51] & B[31];
    assign stage0_r52_c30 = A[52] & B[30];
    assign stage0_r53_c29 = A[53] & B[29];
    assign stage0_r54_c28 = A[54] & B[28];
    assign stage0_r55_c27 = A[55] & B[27];
    assign stage0_r56_c26 = A[56] & B[26];
    assign stage0_r57_c25 = A[57] & B[25];
    assign stage0_r58_c24 = A[58] & B[24];
    assign stage0_r59_c23 = A[59] & B[23];
    assign stage0_r60_c22 = A[60] & B[22];
    assign stage0_r61_c21 = A[61] & B[21];
    assign stage0_r62_c20 = A[62] & B[20];
    assign stage0_r63_c19 = A[63] & B[19];
    assign stage0_r64_c18 = A[64] & B[18];
    assign stage0_r65_c17 = A[65] & B[17];
    assign stage0_r66_c16 = A[66] & B[16];
    assign stage0_r67_c15 = A[67] & B[15];
    assign stage0_r68_c14 = A[68] & B[14];
    assign stage0_r69_c13 = A[69] & B[13];
    assign stage0_r70_c12 = A[70] & B[12];
    assign stage0_r71_c11 = A[71] & B[11];
    assign stage0_r43_c40 = A[43] & B[40];
    assign stage0_r44_c39 = A[44] & B[39];
    assign stage0_r45_c38 = A[45] & B[38];
    assign stage0_r46_c37 = A[46] & B[37];
    assign stage0_r47_c36 = A[47] & B[36];
    assign stage0_r48_c35 = A[48] & B[35];
    assign stage0_r49_c34 = A[49] & B[34];
    assign stage0_r50_c33 = A[50] & B[33];
    assign stage0_r51_c32 = A[51] & B[32];
    assign stage0_r52_c31 = A[52] & B[31];
    assign stage0_r53_c30 = A[53] & B[30];
    assign stage0_r54_c29 = A[54] & B[29];
    assign stage0_r55_c28 = A[55] & B[28];
    assign stage0_r56_c27 = A[56] & B[27];
    assign stage0_r57_c26 = A[57] & B[26];
    assign stage0_r58_c25 = A[58] & B[25];
    assign stage0_r59_c24 = A[59] & B[24];
    assign stage0_r60_c23 = A[60] & B[23];
    assign stage0_r61_c22 = A[61] & B[22];
    assign stage0_r62_c21 = A[62] & B[21];
    assign stage0_r63_c20 = A[63] & B[20];
    assign stage0_r64_c19 = A[64] & B[19];
    assign stage0_r65_c18 = A[65] & B[18];
    assign stage0_r66_c17 = A[66] & B[17];
    assign stage0_r67_c16 = A[67] & B[16];
    assign stage0_r68_c15 = A[68] & B[15];
    assign stage0_r69_c14 = A[69] & B[14];
    assign stage0_r70_c13 = A[70] & B[13];
    assign stage0_r71_c12 = A[71] & B[12];
    assign stage0_r44_c40 = A[44] & B[40];
    assign stage0_r45_c39 = A[45] & B[39];
    assign stage0_r46_c38 = A[46] & B[38];
    assign stage0_r47_c37 = A[47] & B[37];
    assign stage0_r48_c36 = A[48] & B[36];
    assign stage0_r49_c35 = A[49] & B[35];
    assign stage0_r50_c34 = A[50] & B[34];
    assign stage0_r51_c33 = A[51] & B[33];
    assign stage0_r52_c32 = A[52] & B[32];
    assign stage0_r53_c31 = A[53] & B[31];
    assign stage0_r54_c30 = A[54] & B[30];
    assign stage0_r55_c29 = A[55] & B[29];
    assign stage0_r56_c28 = A[56] & B[28];
    assign stage0_r57_c27 = A[57] & B[27];
    assign stage0_r58_c26 = A[58] & B[26];
    assign stage0_r59_c25 = A[59] & B[25];
    assign stage0_r60_c24 = A[60] & B[24];
    assign stage0_r61_c23 = A[61] & B[23];
    assign stage0_r62_c22 = A[62] & B[22];
    assign stage0_r63_c21 = A[63] & B[21];
    assign stage0_r64_c20 = A[64] & B[20];
    assign stage0_r65_c19 = A[65] & B[19];
    assign stage0_r66_c18 = A[66] & B[18];
    assign stage0_r67_c17 = A[67] & B[17];
    assign stage0_r68_c16 = A[68] & B[16];
    assign stage0_r69_c15 = A[69] & B[15];
    assign stage0_r70_c14 = A[70] & B[14];
    assign stage0_r71_c13 = A[71] & B[13];
    assign stage0_r45_c40 = A[45] & B[40];
    assign stage0_r46_c39 = A[46] & B[39];
    assign stage0_r47_c38 = A[47] & B[38];
    assign stage0_r48_c37 = A[48] & B[37];
    assign stage0_r49_c36 = A[49] & B[36];
    assign stage0_r50_c35 = A[50] & B[35];
    assign stage0_r51_c34 = A[51] & B[34];
    assign stage0_r52_c33 = A[52] & B[33];
    assign stage0_r53_c32 = A[53] & B[32];
    assign stage0_r54_c31 = A[54] & B[31];
    assign stage0_r55_c30 = A[55] & B[30];
    assign stage0_r56_c29 = A[56] & B[29];
    assign stage0_r57_c28 = A[57] & B[28];
    assign stage0_r58_c27 = A[58] & B[27];
    assign stage0_r59_c26 = A[59] & B[26];
    assign stage0_r60_c25 = A[60] & B[25];
    assign stage0_r61_c24 = A[61] & B[24];
    assign stage0_r62_c23 = A[62] & B[23];
    assign stage0_r63_c22 = A[63] & B[22];
    assign stage0_r64_c21 = A[64] & B[21];
    assign stage0_r65_c20 = A[65] & B[20];
    assign stage0_r66_c19 = A[66] & B[19];
    assign stage0_r67_c18 = A[67] & B[18];
    assign stage0_r68_c17 = A[68] & B[17];
    assign stage0_r69_c16 = A[69] & B[16];
    assign stage0_r70_c15 = A[70] & B[15];
    assign stage0_r71_c14 = A[71] & B[14];
    assign stage0_r46_c40 = A[46] & B[40];
    assign stage0_r47_c39 = A[47] & B[39];
    assign stage0_r48_c38 = A[48] & B[38];
    assign stage0_r49_c37 = A[49] & B[37];
    assign stage0_r50_c36 = A[50] & B[36];
    assign stage0_r51_c35 = A[51] & B[35];
    assign stage0_r52_c34 = A[52] & B[34];
    assign stage0_r53_c33 = A[53] & B[33];
    assign stage0_r54_c32 = A[54] & B[32];
    assign stage0_r55_c31 = A[55] & B[31];
    assign stage0_r56_c30 = A[56] & B[30];
    assign stage0_r57_c29 = A[57] & B[29];
    assign stage0_r58_c28 = A[58] & B[28];
    assign stage0_r59_c27 = A[59] & B[27];
    assign stage0_r60_c26 = A[60] & B[26];
    assign stage0_r61_c25 = A[61] & B[25];
    assign stage0_r62_c24 = A[62] & B[24];
    assign stage0_r63_c23 = A[63] & B[23];
    assign stage0_r64_c22 = A[64] & B[22];
    assign stage0_r65_c21 = A[65] & B[21];
    assign stage0_r66_c20 = A[66] & B[20];
    assign stage0_r67_c19 = A[67] & B[19];
    assign stage0_r68_c18 = A[68] & B[18];
    assign stage0_r69_c17 = A[69] & B[17];
    assign stage0_r70_c16 = A[70] & B[16];
    assign stage0_r71_c15 = A[71] & B[15];
    assign stage0_r47_c40 = A[47] & B[40];
    assign stage0_r48_c39 = A[48] & B[39];
    assign stage0_r49_c38 = A[49] & B[38];
    assign stage0_r50_c37 = A[50] & B[37];
    assign stage0_r51_c36 = A[51] & B[36];
    assign stage0_r52_c35 = A[52] & B[35];
    assign stage0_r53_c34 = A[53] & B[34];
    assign stage0_r54_c33 = A[54] & B[33];
    assign stage0_r55_c32 = A[55] & B[32];
    assign stage0_r56_c31 = A[56] & B[31];
    assign stage0_r57_c30 = A[57] & B[30];
    assign stage0_r58_c29 = A[58] & B[29];
    assign stage0_r59_c28 = A[59] & B[28];
    assign stage0_r60_c27 = A[60] & B[27];
    assign stage0_r61_c26 = A[61] & B[26];
    assign stage0_r62_c25 = A[62] & B[25];
    assign stage0_r63_c24 = A[63] & B[24];
    assign stage0_r64_c23 = A[64] & B[23];
    assign stage0_r65_c22 = A[65] & B[22];
    assign stage0_r66_c21 = A[66] & B[21];
    assign stage0_r67_c20 = A[67] & B[20];
    assign stage0_r68_c19 = A[68] & B[19];
    assign stage0_r69_c18 = A[69] & B[18];
    assign stage0_r70_c17 = A[70] & B[17];
    assign stage0_r71_c16 = A[71] & B[16];
    assign stage0_r48_c40 = A[48] & B[40];
    assign stage0_r49_c39 = A[49] & B[39];
    assign stage0_r50_c38 = A[50] & B[38];
    assign stage0_r51_c37 = A[51] & B[37];
    assign stage0_r52_c36 = A[52] & B[36];
    assign stage0_r53_c35 = A[53] & B[35];
    assign stage0_r54_c34 = A[54] & B[34];
    assign stage0_r55_c33 = A[55] & B[33];
    assign stage0_r56_c32 = A[56] & B[32];
    assign stage0_r57_c31 = A[57] & B[31];
    assign stage0_r58_c30 = A[58] & B[30];
    assign stage0_r59_c29 = A[59] & B[29];
    assign stage0_r60_c28 = A[60] & B[28];
    assign stage0_r61_c27 = A[61] & B[27];
    assign stage0_r62_c26 = A[62] & B[26];
    assign stage0_r63_c25 = A[63] & B[25];
    assign stage0_r64_c24 = A[64] & B[24];
    assign stage0_r65_c23 = A[65] & B[23];
    assign stage0_r66_c22 = A[66] & B[22];
    assign stage0_r67_c21 = A[67] & B[21];
    assign stage0_r68_c20 = A[68] & B[20];
    assign stage0_r69_c19 = A[69] & B[19];
    assign stage0_r70_c18 = A[70] & B[18];
    assign stage0_r71_c17 = A[71] & B[17];
    assign stage0_r49_c40 = A[49] & B[40];
    assign stage0_r50_c39 = A[50] & B[39];
    assign stage0_r51_c38 = A[51] & B[38];
    assign stage0_r52_c37 = A[52] & B[37];
    assign stage0_r53_c36 = A[53] & B[36];
    assign stage0_r54_c35 = A[54] & B[35];
    assign stage0_r55_c34 = A[55] & B[34];
    assign stage0_r56_c33 = A[56] & B[33];
    assign stage0_r57_c32 = A[57] & B[32];
    assign stage0_r58_c31 = A[58] & B[31];
    assign stage0_r59_c30 = A[59] & B[30];
    assign stage0_r60_c29 = A[60] & B[29];
    assign stage0_r61_c28 = A[61] & B[28];
    assign stage0_r62_c27 = A[62] & B[27];
    assign stage0_r63_c26 = A[63] & B[26];
    assign stage0_r64_c25 = A[64] & B[25];
    assign stage0_r65_c24 = A[65] & B[24];
    assign stage0_r66_c23 = A[66] & B[23];
    assign stage0_r67_c22 = A[67] & B[22];
    assign stage0_r68_c21 = A[68] & B[21];
    assign stage0_r69_c20 = A[69] & B[20];
    assign stage0_r70_c19 = A[70] & B[19];
    assign stage0_r71_c18 = A[71] & B[18];
    assign stage0_r50_c40 = A[50] & B[40];
    assign stage0_r51_c39 = A[51] & B[39];
    assign stage0_r52_c38 = A[52] & B[38];
    assign stage0_r53_c37 = A[53] & B[37];
    assign stage0_r54_c36 = A[54] & B[36];
    assign stage0_r55_c35 = A[55] & B[35];
    assign stage0_r56_c34 = A[56] & B[34];
    assign stage0_r57_c33 = A[57] & B[33];
    assign stage0_r58_c32 = A[58] & B[32];
    assign stage0_r59_c31 = A[59] & B[31];
    assign stage0_r60_c30 = A[60] & B[30];
    assign stage0_r61_c29 = A[61] & B[29];
    assign stage0_r62_c28 = A[62] & B[28];
    assign stage0_r63_c27 = A[63] & B[27];
    assign stage0_r64_c26 = A[64] & B[26];
    assign stage0_r65_c25 = A[65] & B[25];
    assign stage0_r66_c24 = A[66] & B[24];
    assign stage0_r67_c23 = A[67] & B[23];
    assign stage0_r68_c22 = A[68] & B[22];
    assign stage0_r69_c21 = A[69] & B[21];
    assign stage0_r70_c20 = A[70] & B[20];
    assign stage0_r71_c19 = A[71] & B[19];
    assign stage0_r51_c40 = A[51] & B[40];
    assign stage0_r52_c39 = A[52] & B[39];
    assign stage0_r53_c38 = A[53] & B[38];
    assign stage0_r54_c37 = A[54] & B[37];
    assign stage0_r55_c36 = A[55] & B[36];
    assign stage0_r56_c35 = A[56] & B[35];
    assign stage0_r57_c34 = A[57] & B[34];
    assign stage0_r58_c33 = A[58] & B[33];
    assign stage0_r59_c32 = A[59] & B[32];
    assign stage0_r60_c31 = A[60] & B[31];
    assign stage0_r61_c30 = A[61] & B[30];
    assign stage0_r62_c29 = A[62] & B[29];
    assign stage0_r63_c28 = A[63] & B[28];
    assign stage0_r64_c27 = A[64] & B[27];
    assign stage0_r65_c26 = A[65] & B[26];
    assign stage0_r66_c25 = A[66] & B[25];
    assign stage0_r67_c24 = A[67] & B[24];
    assign stage0_r68_c23 = A[68] & B[23];
    assign stage0_r69_c22 = A[69] & B[22];
    assign stage0_r70_c21 = A[70] & B[21];
    assign stage0_r71_c20 = A[71] & B[20];
    assign stage0_r52_c40 = A[52] & B[40];
    assign stage0_r53_c39 = A[53] & B[39];
    assign stage0_r54_c38 = A[54] & B[38];
    assign stage0_r55_c37 = A[55] & B[37];
    assign stage0_r56_c36 = A[56] & B[36];
    assign stage0_r57_c35 = A[57] & B[35];
    assign stage0_r58_c34 = A[58] & B[34];
    assign stage0_r59_c33 = A[59] & B[33];
    assign stage0_r60_c32 = A[60] & B[32];
    assign stage0_r61_c31 = A[61] & B[31];
    assign stage0_r62_c30 = A[62] & B[30];
    assign stage0_r63_c29 = A[63] & B[29];
    assign stage0_r64_c28 = A[64] & B[28];
    assign stage0_r65_c27 = A[65] & B[27];
    assign stage0_r66_c26 = A[66] & B[26];
    assign stage0_r67_c25 = A[67] & B[25];
    assign stage0_r68_c24 = A[68] & B[24];
    assign stage0_r69_c23 = A[69] & B[23];
    assign stage0_r70_c22 = A[70] & B[22];
    assign stage0_r71_c21 = A[71] & B[21];
    assign stage0_r53_c40 = A[53] & B[40];
    assign stage0_r54_c39 = A[54] & B[39];
    assign stage0_r55_c38 = A[55] & B[38];
    assign stage0_r56_c37 = A[56] & B[37];
    assign stage0_r57_c36 = A[57] & B[36];
    assign stage0_r58_c35 = A[58] & B[35];
    assign stage0_r59_c34 = A[59] & B[34];
    assign stage0_r60_c33 = A[60] & B[33];
    assign stage0_r61_c32 = A[61] & B[32];
    assign stage0_r62_c31 = A[62] & B[31];
    assign stage0_r63_c30 = A[63] & B[30];
    assign stage0_r64_c29 = A[64] & B[29];
    assign stage0_r65_c28 = A[65] & B[28];
    assign stage0_r66_c27 = A[66] & B[27];
    assign stage0_r67_c26 = A[67] & B[26];
    assign stage0_r68_c25 = A[68] & B[25];
    assign stage0_r69_c24 = A[69] & B[24];
    assign stage0_r70_c23 = A[70] & B[23];
    assign stage0_r71_c22 = A[71] & B[22];
    assign stage0_r54_c40 = A[54] & B[40];
    assign stage0_r55_c39 = A[55] & B[39];
    assign stage0_r56_c38 = A[56] & B[38];
    assign stage0_r57_c37 = A[57] & B[37];
    assign stage0_r58_c36 = A[58] & B[36];
    assign stage0_r59_c35 = A[59] & B[35];
    assign stage0_r60_c34 = A[60] & B[34];
    assign stage0_r61_c33 = A[61] & B[33];
    assign stage0_r62_c32 = A[62] & B[32];
    assign stage0_r63_c31 = A[63] & B[31];
    assign stage0_r64_c30 = A[64] & B[30];
    assign stage0_r65_c29 = A[65] & B[29];
    assign stage0_r66_c28 = A[66] & B[28];
    assign stage0_r67_c27 = A[67] & B[27];
    assign stage0_r68_c26 = A[68] & B[26];
    assign stage0_r69_c25 = A[69] & B[25];
    assign stage0_r70_c24 = A[70] & B[24];
    assign stage0_r71_c23 = A[71] & B[23];
    assign stage0_r55_c40 = A[55] & B[40];
    assign stage0_r56_c39 = A[56] & B[39];
    assign stage0_r57_c38 = A[57] & B[38];
    assign stage0_r58_c37 = A[58] & B[37];
    assign stage0_r59_c36 = A[59] & B[36];
    assign stage0_r60_c35 = A[60] & B[35];
    assign stage0_r61_c34 = A[61] & B[34];
    assign stage0_r62_c33 = A[62] & B[33];
    assign stage0_r63_c32 = A[63] & B[32];
    assign stage0_r64_c31 = A[64] & B[31];
    assign stage0_r65_c30 = A[65] & B[30];
    assign stage0_r66_c29 = A[66] & B[29];
    assign stage0_r67_c28 = A[67] & B[28];
    assign stage0_r68_c27 = A[68] & B[27];
    assign stage0_r69_c26 = A[69] & B[26];
    assign stage0_r70_c25 = A[70] & B[25];
    assign stage0_r71_c24 = A[71] & B[24];
    assign stage0_r56_c40 = A[56] & B[40];
    assign stage0_r57_c39 = A[57] & B[39];
    assign stage0_r58_c38 = A[58] & B[38];
    assign stage0_r59_c37 = A[59] & B[37];
    assign stage0_r60_c36 = A[60] & B[36];
    assign stage0_r61_c35 = A[61] & B[35];
    assign stage0_r62_c34 = A[62] & B[34];
    assign stage0_r63_c33 = A[63] & B[33];
    assign stage0_r64_c32 = A[64] & B[32];
    assign stage0_r65_c31 = A[65] & B[31];
    assign stage0_r66_c30 = A[66] & B[30];
    assign stage0_r67_c29 = A[67] & B[29];
    assign stage0_r68_c28 = A[68] & B[28];
    assign stage0_r69_c27 = A[69] & B[27];
    assign stage0_r70_c26 = A[70] & B[26];
    assign stage0_r71_c25 = A[71] & B[25];
    assign stage0_r57_c40 = A[57] & B[40];
    assign stage0_r58_c39 = A[58] & B[39];
    assign stage0_r59_c38 = A[59] & B[38];
    assign stage0_r60_c37 = A[60] & B[37];
    assign stage0_r61_c36 = A[61] & B[36];
    assign stage0_r62_c35 = A[62] & B[35];
    assign stage0_r63_c34 = A[63] & B[34];
    assign stage0_r64_c33 = A[64] & B[33];
    assign stage0_r65_c32 = A[65] & B[32];
    assign stage0_r66_c31 = A[66] & B[31];
    assign stage0_r67_c30 = A[67] & B[30];
    assign stage0_r68_c29 = A[68] & B[29];
    assign stage0_r69_c28 = A[69] & B[28];
    assign stage0_r70_c27 = A[70] & B[27];
    assign stage0_r71_c26 = A[71] & B[26];
    assign stage0_r58_c40 = A[58] & B[40];
    assign stage0_r59_c39 = A[59] & B[39];
    assign stage0_r60_c38 = A[60] & B[38];
    assign stage0_r61_c37 = A[61] & B[37];
    assign stage0_r62_c36 = A[62] & B[36];
    assign stage0_r63_c35 = A[63] & B[35];
    assign stage0_r64_c34 = A[64] & B[34];
    assign stage0_r65_c33 = A[65] & B[33];
    assign stage0_r66_c32 = A[66] & B[32];
    assign stage0_r67_c31 = A[67] & B[31];
    assign stage0_r68_c30 = A[68] & B[30];
    assign stage0_r69_c29 = A[69] & B[29];
    assign stage0_r70_c28 = A[70] & B[28];
    assign stage0_r71_c27 = A[71] & B[27];
    assign stage0_r59_c40 = A[59] & B[40];
    assign stage0_r60_c39 = A[60] & B[39];
    assign stage0_r61_c38 = A[61] & B[38];
    assign stage0_r62_c37 = A[62] & B[37];
    assign stage0_r63_c36 = A[63] & B[36];
    assign stage0_r64_c35 = A[64] & B[35];
    assign stage0_r65_c34 = A[65] & B[34];
    assign stage0_r66_c33 = A[66] & B[33];
    assign stage0_r67_c32 = A[67] & B[32];
    assign stage0_r68_c31 = A[68] & B[31];
    assign stage0_r69_c30 = A[69] & B[30];
    assign stage0_r70_c29 = A[70] & B[29];
    assign stage0_r71_c28 = A[71] & B[28];
    assign stage0_r60_c40 = A[60] & B[40];
    assign stage0_r61_c39 = A[61] & B[39];
    assign stage0_r62_c38 = A[62] & B[38];
    assign stage0_r63_c37 = A[63] & B[37];
    assign stage0_r64_c36 = A[64] & B[36];
    assign stage0_r65_c35 = A[65] & B[35];
    assign stage0_r66_c34 = A[66] & B[34];
    assign stage0_r67_c33 = A[67] & B[33];
    assign stage0_r68_c32 = A[68] & B[32];
    assign stage0_r69_c31 = A[69] & B[31];
    assign stage0_r70_c30 = A[70] & B[30];
    assign stage0_r71_c29 = A[71] & B[29];
    assign stage0_r61_c40 = A[61] & B[40];
    assign stage0_r62_c39 = A[62] & B[39];
    assign stage0_r63_c38 = A[63] & B[38];
    assign stage0_r64_c37 = A[64] & B[37];
    assign stage0_r65_c36 = A[65] & B[36];
    assign stage0_r66_c35 = A[66] & B[35];
    assign stage0_r67_c34 = A[67] & B[34];
    assign stage0_r68_c33 = A[68] & B[33];
    assign stage0_r69_c32 = A[69] & B[32];
    assign stage0_r70_c31 = A[70] & B[31];
    assign stage0_r71_c30 = A[71] & B[30];
    assign stage0_r62_c40 = A[62] & B[40];
    assign stage0_r63_c39 = A[63] & B[39];
    assign stage0_r64_c38 = A[64] & B[38];
    assign stage0_r65_c37 = A[65] & B[37];
    assign stage0_r66_c36 = A[66] & B[36];
    assign stage0_r67_c35 = A[67] & B[35];
    assign stage0_r68_c34 = A[68] & B[34];
    assign stage0_r69_c33 = A[69] & B[33];
    assign stage0_r70_c32 = A[70] & B[32];
    assign stage0_r71_c31 = A[71] & B[31];
    assign stage0_r63_c40 = A[63] & B[40];
    assign stage0_r64_c39 = A[64] & B[39];
    assign stage0_r65_c38 = A[65] & B[38];
    assign stage0_r66_c37 = A[66] & B[37];
    assign stage0_r67_c36 = A[67] & B[36];
    assign stage0_r68_c35 = A[68] & B[35];
    assign stage0_r69_c34 = A[69] & B[34];
    assign stage0_r70_c33 = A[70] & B[33];
    assign stage0_r71_c32 = A[71] & B[32];
    assign stage0_r64_c40 = A[64] & B[40];
    assign stage0_r65_c39 = A[65] & B[39];
    assign stage0_r66_c38 = A[66] & B[38];
    assign stage0_r67_c37 = A[67] & B[37];
    assign stage0_r68_c36 = A[68] & B[36];
    assign stage0_r69_c35 = A[69] & B[35];
    assign stage0_r70_c34 = A[70] & B[34];
    assign stage0_r71_c33 = A[71] & B[33];
    assign stage0_r65_c40 = A[65] & B[40];
    assign stage0_r66_c39 = A[66] & B[39];
    assign stage0_r67_c38 = A[67] & B[38];
    assign stage0_r68_c37 = A[68] & B[37];
    assign stage0_r69_c36 = A[69] & B[36];
    assign stage0_r70_c35 = A[70] & B[35];
    assign stage0_r71_c34 = A[71] & B[34];
    assign stage0_r66_c40 = A[66] & B[40];
    assign stage0_r67_c39 = A[67] & B[39];
    assign stage0_r68_c38 = A[68] & B[38];
    assign stage0_r69_c37 = A[69] & B[37];
    assign stage0_r70_c36 = A[70] & B[36];
    assign stage0_r71_c35 = A[71] & B[35];
    assign stage0_r67_c40 = A[67] & B[40];
    assign stage0_r68_c39 = A[68] & B[39];
    assign stage0_r69_c38 = A[69] & B[38];
    assign stage0_r70_c37 = A[70] & B[37];
    assign stage0_r71_c36 = A[71] & B[36];
    assign stage0_r68_c40 = A[68] & B[40];
    assign stage0_r69_c39 = A[69] & B[39];
    assign stage0_r70_c38 = A[70] & B[38];
    assign stage0_r71_c37 = A[71] & B[37];
    assign stage0_r69_c40 = A[69] & B[40];
    assign stage0_r70_c39 = A[70] & B[39];
    assign stage0_r71_c38 = A[71] & B[38];
    assign stage0_r70_c40 = A[70] & B[40];
    assign stage0_r71_c39 = A[71] & B[39];
    assign stage0_r71_c40 = A[71] & B[40];
    HA ha_0(.A(stage0_r0_c1), .B(stage0_r1_c0), .So(stage1_c1_s_ha0), .Co(stage1_c1_c_ha0));
    FA fa_0(.A(stage0_r0_c2), .B(stage0_r1_c1), .C(stage0_r2_c0), .So(stage1_c2_s_fa0), .Co(stage1_c2_c_fa0));
    FA fa_1(.A(stage0_r0_c3), .B(stage0_r1_c2), .C(stage0_r2_c1), .So(stage1_c3_s_fa0), .Co(stage1_c3_c_fa0));
    FA fa_2(.A(stage0_r0_c4), .B(stage0_r1_c3), .C(stage0_r2_c2), .So(stage1_c4_s_fa0), .Co(stage1_c4_c_fa0));
    HA ha_1(.A(stage0_r3_c1), .B(stage0_r4_c0), .So(stage1_c4_s_ha0), .Co(stage1_c4_c_ha0));
    FA fa_3(.A(stage0_r0_c5), .B(stage0_r1_c4), .C(stage0_r2_c3), .So(stage1_c5_s_fa0), .Co(stage1_c5_c_fa0));
    FA fa_4(.A(stage0_r3_c2), .B(stage0_r4_c1), .C(stage0_r5_c0), .So(stage1_c5_s_fa1), .Co(stage1_c5_c_fa1));
    FA fa_5(.A(stage0_r0_c6), .B(stage0_r1_c5), .C(stage0_r2_c4), .So(stage1_c6_s_fa0), .Co(stage1_c6_c_fa0));
    FA fa_6(.A(stage0_r3_c3), .B(stage0_r4_c2), .C(stage0_r5_c1), .So(stage1_c6_s_fa1), .Co(stage1_c6_c_fa1));
    FA fa_7(.A(stage0_r0_c7), .B(stage0_r1_c6), .C(stage0_r2_c5), .So(stage1_c7_s_fa0), .Co(stage1_c7_c_fa0));
    FA fa_8(.A(stage0_r3_c4), .B(stage0_r4_c3), .C(stage0_r5_c2), .So(stage1_c7_s_fa1), .Co(stage1_c7_c_fa1));
    HA ha_2(.A(stage0_r6_c1), .B(stage0_r7_c0), .So(stage1_c7_s_ha0), .Co(stage1_c7_c_ha0));
    FA fa_9(.A(stage0_r0_c8), .B(stage0_r1_c7), .C(stage0_r2_c6), .So(stage1_c8_s_fa0), .Co(stage1_c8_c_fa0));
    FA fa_10(.A(stage0_r3_c5), .B(stage0_r4_c4), .C(stage0_r5_c3), .So(stage1_c8_s_fa1), .Co(stage1_c8_c_fa1));
    FA fa_11(.A(stage0_r6_c2), .B(stage0_r7_c1), .C(stage0_r8_c0), .So(stage1_c8_s_fa2), .Co(stage1_c8_c_fa2));
    FA fa_12(.A(stage0_r0_c9), .B(stage0_r1_c8), .C(stage0_r2_c7), .So(stage1_c9_s_fa0), .Co(stage1_c9_c_fa0));
    FA fa_13(.A(stage0_r3_c6), .B(stage0_r4_c5), .C(stage0_r5_c4), .So(stage1_c9_s_fa1), .Co(stage1_c9_c_fa1));
    FA fa_14(.A(stage0_r6_c3), .B(stage0_r7_c2), .C(stage0_r8_c1), .So(stage1_c9_s_fa2), .Co(stage1_c9_c_fa2));
    FA fa_15(.A(stage0_r0_c10), .B(stage0_r1_c9), .C(stage0_r2_c8), .So(stage1_c10_s_fa0), .Co(stage1_c10_c_fa0));
    FA fa_16(.A(stage0_r3_c7), .B(stage0_r4_c6), .C(stage0_r5_c5), .So(stage1_c10_s_fa1), .Co(stage1_c10_c_fa1));
    FA fa_17(.A(stage0_r6_c4), .B(stage0_r7_c3), .C(stage0_r8_c2), .So(stage1_c10_s_fa2), .Co(stage1_c10_c_fa2));
    HA ha_3(.A(stage0_r9_c1), .B(stage0_r10_c0), .So(stage1_c10_s_ha0), .Co(stage1_c10_c_ha0));
    FA fa_18(.A(stage0_r0_c11), .B(stage0_r1_c10), .C(stage0_r2_c9), .So(stage1_c11_s_fa0), .Co(stage1_c11_c_fa0));
    FA fa_19(.A(stage0_r3_c8), .B(stage0_r4_c7), .C(stage0_r5_c6), .So(stage1_c11_s_fa1), .Co(stage1_c11_c_fa1));
    FA fa_20(.A(stage0_r6_c5), .B(stage0_r7_c4), .C(stage0_r8_c3), .So(stage1_c11_s_fa2), .Co(stage1_c11_c_fa2));
    FA fa_21(.A(stage0_r9_c2), .B(stage0_r10_c1), .C(stage0_r11_c0), .So(stage1_c11_s_fa3), .Co(stage1_c11_c_fa3));
    FA fa_22(.A(stage0_r0_c12), .B(stage0_r1_c11), .C(stage0_r2_c10), .So(stage1_c12_s_fa0), .Co(stage1_c12_c_fa0));
    FA fa_23(.A(stage0_r3_c9), .B(stage0_r4_c8), .C(stage0_r5_c7), .So(stage1_c12_s_fa1), .Co(stage1_c12_c_fa1));
    FA fa_24(.A(stage0_r6_c6), .B(stage0_r7_c5), .C(stage0_r8_c4), .So(stage1_c12_s_fa2), .Co(stage1_c12_c_fa2));
    FA fa_25(.A(stage0_r9_c3), .B(stage0_r10_c2), .C(stage0_r11_c1), .So(stage1_c12_s_fa3), .Co(stage1_c12_c_fa3));
    FA fa_26(.A(stage0_r0_c13), .B(stage0_r1_c12), .C(stage0_r2_c11), .So(stage1_c13_s_fa0), .Co(stage1_c13_c_fa0));
    FA fa_27(.A(stage0_r3_c10), .B(stage0_r4_c9), .C(stage0_r5_c8), .So(stage1_c13_s_fa1), .Co(stage1_c13_c_fa1));
    FA fa_28(.A(stage0_r6_c7), .B(stage0_r7_c6), .C(stage0_r8_c5), .So(stage1_c13_s_fa2), .Co(stage1_c13_c_fa2));
    FA fa_29(.A(stage0_r9_c4), .B(stage0_r10_c3), .C(stage0_r11_c2), .So(stage1_c13_s_fa3), .Co(stage1_c13_c_fa3));
    HA ha_4(.A(stage0_r12_c1), .B(stage0_r13_c0), .So(stage1_c13_s_ha0), .Co(stage1_c13_c_ha0));
    FA fa_30(.A(stage0_r0_c14), .B(stage0_r1_c13), .C(stage0_r2_c12), .So(stage1_c14_s_fa0), .Co(stage1_c14_c_fa0));
    FA fa_31(.A(stage0_r3_c11), .B(stage0_r4_c10), .C(stage0_r5_c9), .So(stage1_c14_s_fa1), .Co(stage1_c14_c_fa1));
    FA fa_32(.A(stage0_r6_c8), .B(stage0_r7_c7), .C(stage0_r8_c6), .So(stage1_c14_s_fa2), .Co(stage1_c14_c_fa2));
    FA fa_33(.A(stage0_r9_c5), .B(stage0_r10_c4), .C(stage0_r11_c3), .So(stage1_c14_s_fa3), .Co(stage1_c14_c_fa3));
    FA fa_34(.A(stage0_r12_c2), .B(stage0_r13_c1), .C(stage0_r14_c0), .So(stage1_c14_s_fa4), .Co(stage1_c14_c_fa4));
    FA fa_35(.A(stage0_r0_c15), .B(stage0_r1_c14), .C(stage0_r2_c13), .So(stage1_c15_s_fa0), .Co(stage1_c15_c_fa0));
    FA fa_36(.A(stage0_r3_c12), .B(stage0_r4_c11), .C(stage0_r5_c10), .So(stage1_c15_s_fa1), .Co(stage1_c15_c_fa1));
    FA fa_37(.A(stage0_r6_c9), .B(stage0_r7_c8), .C(stage0_r8_c7), .So(stage1_c15_s_fa2), .Co(stage1_c15_c_fa2));
    FA fa_38(.A(stage0_r9_c6), .B(stage0_r10_c5), .C(stage0_r11_c4), .So(stage1_c15_s_fa3), .Co(stage1_c15_c_fa3));
    FA fa_39(.A(stage0_r12_c3), .B(stage0_r13_c2), .C(stage0_r14_c1), .So(stage1_c15_s_fa4), .Co(stage1_c15_c_fa4));
    FA fa_40(.A(stage0_r0_c16), .B(stage0_r1_c15), .C(stage0_r2_c14), .So(stage1_c16_s_fa0), .Co(stage1_c16_c_fa0));
    FA fa_41(.A(stage0_r3_c13), .B(stage0_r4_c12), .C(stage0_r5_c11), .So(stage1_c16_s_fa1), .Co(stage1_c16_c_fa1));
    FA fa_42(.A(stage0_r6_c10), .B(stage0_r7_c9), .C(stage0_r8_c8), .So(stage1_c16_s_fa2), .Co(stage1_c16_c_fa2));
    FA fa_43(.A(stage0_r9_c7), .B(stage0_r10_c6), .C(stage0_r11_c5), .So(stage1_c16_s_fa3), .Co(stage1_c16_c_fa3));
    FA fa_44(.A(stage0_r12_c4), .B(stage0_r13_c3), .C(stage0_r14_c2), .So(stage1_c16_s_fa4), .Co(stage1_c16_c_fa4));
    HA ha_5(.A(stage0_r15_c1), .B(stage0_r16_c0), .So(stage1_c16_s_ha0), .Co(stage1_c16_c_ha0));
    FA fa_45(.A(stage0_r0_c17), .B(stage0_r1_c16), .C(stage0_r2_c15), .So(stage1_c17_s_fa0), .Co(stage1_c17_c_fa0));
    FA fa_46(.A(stage0_r3_c14), .B(stage0_r4_c13), .C(stage0_r5_c12), .So(stage1_c17_s_fa1), .Co(stage1_c17_c_fa1));
    FA fa_47(.A(stage0_r6_c11), .B(stage0_r7_c10), .C(stage0_r8_c9), .So(stage1_c17_s_fa2), .Co(stage1_c17_c_fa2));
    FA fa_48(.A(stage0_r9_c8), .B(stage0_r10_c7), .C(stage0_r11_c6), .So(stage1_c17_s_fa3), .Co(stage1_c17_c_fa3));
    FA fa_49(.A(stage0_r12_c5), .B(stage0_r13_c4), .C(stage0_r14_c3), .So(stage1_c17_s_fa4), .Co(stage1_c17_c_fa4));
    FA fa_50(.A(stage0_r15_c2), .B(stage0_r16_c1), .C(stage0_r17_c0), .So(stage1_c17_s_fa5), .Co(stage1_c17_c_fa5));
    FA fa_51(.A(stage0_r0_c18), .B(stage0_r1_c17), .C(stage0_r2_c16), .So(stage1_c18_s_fa0), .Co(stage1_c18_c_fa0));
    FA fa_52(.A(stage0_r3_c15), .B(stage0_r4_c14), .C(stage0_r5_c13), .So(stage1_c18_s_fa1), .Co(stage1_c18_c_fa1));
    FA fa_53(.A(stage0_r6_c12), .B(stage0_r7_c11), .C(stage0_r8_c10), .So(stage1_c18_s_fa2), .Co(stage1_c18_c_fa2));
    FA fa_54(.A(stage0_r9_c9), .B(stage0_r10_c8), .C(stage0_r11_c7), .So(stage1_c18_s_fa3), .Co(stage1_c18_c_fa3));
    FA fa_55(.A(stage0_r12_c6), .B(stage0_r13_c5), .C(stage0_r14_c4), .So(stage1_c18_s_fa4), .Co(stage1_c18_c_fa4));
    FA fa_56(.A(stage0_r15_c3), .B(stage0_r16_c2), .C(stage0_r17_c1), .So(stage1_c18_s_fa5), .Co(stage1_c18_c_fa5));
    FA fa_57(.A(stage0_r0_c19), .B(stage0_r1_c18), .C(stage0_r2_c17), .So(stage1_c19_s_fa0), .Co(stage1_c19_c_fa0));
    FA fa_58(.A(stage0_r3_c16), .B(stage0_r4_c15), .C(stage0_r5_c14), .So(stage1_c19_s_fa1), .Co(stage1_c19_c_fa1));
    FA fa_59(.A(stage0_r6_c13), .B(stage0_r7_c12), .C(stage0_r8_c11), .So(stage1_c19_s_fa2), .Co(stage1_c19_c_fa2));
    FA fa_60(.A(stage0_r9_c10), .B(stage0_r10_c9), .C(stage0_r11_c8), .So(stage1_c19_s_fa3), .Co(stage1_c19_c_fa3));
    FA fa_61(.A(stage0_r12_c7), .B(stage0_r13_c6), .C(stage0_r14_c5), .So(stage1_c19_s_fa4), .Co(stage1_c19_c_fa4));
    FA fa_62(.A(stage0_r15_c4), .B(stage0_r16_c3), .C(stage0_r17_c2), .So(stage1_c19_s_fa5), .Co(stage1_c19_c_fa5));
    HA ha_6(.A(stage0_r18_c1), .B(stage0_r19_c0), .So(stage1_c19_s_ha0), .Co(stage1_c19_c_ha0));
    FA fa_63(.A(stage0_r0_c20), .B(stage0_r1_c19), .C(stage0_r2_c18), .So(stage1_c20_s_fa0), .Co(stage1_c20_c_fa0));
    FA fa_64(.A(stage0_r3_c17), .B(stage0_r4_c16), .C(stage0_r5_c15), .So(stage1_c20_s_fa1), .Co(stage1_c20_c_fa1));
    FA fa_65(.A(stage0_r6_c14), .B(stage0_r7_c13), .C(stage0_r8_c12), .So(stage1_c20_s_fa2), .Co(stage1_c20_c_fa2));
    FA fa_66(.A(stage0_r9_c11), .B(stage0_r10_c10), .C(stage0_r11_c9), .So(stage1_c20_s_fa3), .Co(stage1_c20_c_fa3));
    FA fa_67(.A(stage0_r12_c8), .B(stage0_r13_c7), .C(stage0_r14_c6), .So(stage1_c20_s_fa4), .Co(stage1_c20_c_fa4));
    FA fa_68(.A(stage0_r15_c5), .B(stage0_r16_c4), .C(stage0_r17_c3), .So(stage1_c20_s_fa5), .Co(stage1_c20_c_fa5));
    FA fa_69(.A(stage0_r18_c2), .B(stage0_r19_c1), .C(stage0_r20_c0), .So(stage1_c20_s_fa6), .Co(stage1_c20_c_fa6));
    FA fa_70(.A(stage0_r0_c21), .B(stage0_r1_c20), .C(stage0_r2_c19), .So(stage1_c21_s_fa0), .Co(stage1_c21_c_fa0));
    FA fa_71(.A(stage0_r3_c18), .B(stage0_r4_c17), .C(stage0_r5_c16), .So(stage1_c21_s_fa1), .Co(stage1_c21_c_fa1));
    FA fa_72(.A(stage0_r6_c15), .B(stage0_r7_c14), .C(stage0_r8_c13), .So(stage1_c21_s_fa2), .Co(stage1_c21_c_fa2));
    FA fa_73(.A(stage0_r9_c12), .B(stage0_r10_c11), .C(stage0_r11_c10), .So(stage1_c21_s_fa3), .Co(stage1_c21_c_fa3));
    FA fa_74(.A(stage0_r12_c9), .B(stage0_r13_c8), .C(stage0_r14_c7), .So(stage1_c21_s_fa4), .Co(stage1_c21_c_fa4));
    FA fa_75(.A(stage0_r15_c6), .B(stage0_r16_c5), .C(stage0_r17_c4), .So(stage1_c21_s_fa5), .Co(stage1_c21_c_fa5));
    FA fa_76(.A(stage0_r18_c3), .B(stage0_r19_c2), .C(stage0_r20_c1), .So(stage1_c21_s_fa6), .Co(stage1_c21_c_fa6));
    FA fa_77(.A(stage0_r0_c22), .B(stage0_r1_c21), .C(stage0_r2_c20), .So(stage1_c22_s_fa0), .Co(stage1_c22_c_fa0));
    FA fa_78(.A(stage0_r3_c19), .B(stage0_r4_c18), .C(stage0_r5_c17), .So(stage1_c22_s_fa1), .Co(stage1_c22_c_fa1));
    FA fa_79(.A(stage0_r6_c16), .B(stage0_r7_c15), .C(stage0_r8_c14), .So(stage1_c22_s_fa2), .Co(stage1_c22_c_fa2));
    FA fa_80(.A(stage0_r9_c13), .B(stage0_r10_c12), .C(stage0_r11_c11), .So(stage1_c22_s_fa3), .Co(stage1_c22_c_fa3));
    FA fa_81(.A(stage0_r12_c10), .B(stage0_r13_c9), .C(stage0_r14_c8), .So(stage1_c22_s_fa4), .Co(stage1_c22_c_fa4));
    FA fa_82(.A(stage0_r15_c7), .B(stage0_r16_c6), .C(stage0_r17_c5), .So(stage1_c22_s_fa5), .Co(stage1_c22_c_fa5));
    FA fa_83(.A(stage0_r18_c4), .B(stage0_r19_c3), .C(stage0_r20_c2), .So(stage1_c22_s_fa6), .Co(stage1_c22_c_fa6));
    HA ha_7(.A(stage0_r21_c1), .B(stage0_r22_c0), .So(stage1_c22_s_ha0), .Co(stage1_c22_c_ha0));
    FA fa_84(.A(stage0_r0_c23), .B(stage0_r1_c22), .C(stage0_r2_c21), .So(stage1_c23_s_fa0), .Co(stage1_c23_c_fa0));
    FA fa_85(.A(stage0_r3_c20), .B(stage0_r4_c19), .C(stage0_r5_c18), .So(stage1_c23_s_fa1), .Co(stage1_c23_c_fa1));
    FA fa_86(.A(stage0_r6_c17), .B(stage0_r7_c16), .C(stage0_r8_c15), .So(stage1_c23_s_fa2), .Co(stage1_c23_c_fa2));
    FA fa_87(.A(stage0_r9_c14), .B(stage0_r10_c13), .C(stage0_r11_c12), .So(stage1_c23_s_fa3), .Co(stage1_c23_c_fa3));
    FA fa_88(.A(stage0_r12_c11), .B(stage0_r13_c10), .C(stage0_r14_c9), .So(stage1_c23_s_fa4), .Co(stage1_c23_c_fa4));
    FA fa_89(.A(stage0_r15_c8), .B(stage0_r16_c7), .C(stage0_r17_c6), .So(stage1_c23_s_fa5), .Co(stage1_c23_c_fa5));
    FA fa_90(.A(stage0_r18_c5), .B(stage0_r19_c4), .C(stage0_r20_c3), .So(stage1_c23_s_fa6), .Co(stage1_c23_c_fa6));
    FA fa_91(.A(stage0_r21_c2), .B(stage0_r22_c1), .C(stage0_r23_c0), .So(stage1_c23_s_fa7), .Co(stage1_c23_c_fa7));
    FA fa_92(.A(stage0_r0_c24), .B(stage0_r1_c23), .C(stage0_r2_c22), .So(stage1_c24_s_fa0), .Co(stage1_c24_c_fa0));
    FA fa_93(.A(stage0_r3_c21), .B(stage0_r4_c20), .C(stage0_r5_c19), .So(stage1_c24_s_fa1), .Co(stage1_c24_c_fa1));
    FA fa_94(.A(stage0_r6_c18), .B(stage0_r7_c17), .C(stage0_r8_c16), .So(stage1_c24_s_fa2), .Co(stage1_c24_c_fa2));
    FA fa_95(.A(stage0_r9_c15), .B(stage0_r10_c14), .C(stage0_r11_c13), .So(stage1_c24_s_fa3), .Co(stage1_c24_c_fa3));
    FA fa_96(.A(stage0_r12_c12), .B(stage0_r13_c11), .C(stage0_r14_c10), .So(stage1_c24_s_fa4), .Co(stage1_c24_c_fa4));
    FA fa_97(.A(stage0_r15_c9), .B(stage0_r16_c8), .C(stage0_r17_c7), .So(stage1_c24_s_fa5), .Co(stage1_c24_c_fa5));
    FA fa_98(.A(stage0_r18_c6), .B(stage0_r19_c5), .C(stage0_r20_c4), .So(stage1_c24_s_fa6), .Co(stage1_c24_c_fa6));
    FA fa_99(.A(stage0_r21_c3), .B(stage0_r22_c2), .C(stage0_r23_c1), .So(stage1_c24_s_fa7), .Co(stage1_c24_c_fa7));
    FA fa_100(.A(stage0_r0_c25), .B(stage0_r1_c24), .C(stage0_r2_c23), .So(stage1_c25_s_fa0), .Co(stage1_c25_c_fa0));
    FA fa_101(.A(stage0_r3_c22), .B(stage0_r4_c21), .C(stage0_r5_c20), .So(stage1_c25_s_fa1), .Co(stage1_c25_c_fa1));
    FA fa_102(.A(stage0_r6_c19), .B(stage0_r7_c18), .C(stage0_r8_c17), .So(stage1_c25_s_fa2), .Co(stage1_c25_c_fa2));
    FA fa_103(.A(stage0_r9_c16), .B(stage0_r10_c15), .C(stage0_r11_c14), .So(stage1_c25_s_fa3), .Co(stage1_c25_c_fa3));
    FA fa_104(.A(stage0_r12_c13), .B(stage0_r13_c12), .C(stage0_r14_c11), .So(stage1_c25_s_fa4), .Co(stage1_c25_c_fa4));
    FA fa_105(.A(stage0_r15_c10), .B(stage0_r16_c9), .C(stage0_r17_c8), .So(stage1_c25_s_fa5), .Co(stage1_c25_c_fa5));
    FA fa_106(.A(stage0_r18_c7), .B(stage0_r19_c6), .C(stage0_r20_c5), .So(stage1_c25_s_fa6), .Co(stage1_c25_c_fa6));
    FA fa_107(.A(stage0_r21_c4), .B(stage0_r22_c3), .C(stage0_r23_c2), .So(stage1_c25_s_fa7), .Co(stage1_c25_c_fa7));
    HA ha_8(.A(stage0_r24_c1), .B(stage0_r25_c0), .So(stage1_c25_s_ha0), .Co(stage1_c25_c_ha0));
    FA fa_108(.A(stage0_r0_c26), .B(stage0_r1_c25), .C(stage0_r2_c24), .So(stage1_c26_s_fa0), .Co(stage1_c26_c_fa0));
    FA fa_109(.A(stage0_r3_c23), .B(stage0_r4_c22), .C(stage0_r5_c21), .So(stage1_c26_s_fa1), .Co(stage1_c26_c_fa1));
    FA fa_110(.A(stage0_r6_c20), .B(stage0_r7_c19), .C(stage0_r8_c18), .So(stage1_c26_s_fa2), .Co(stage1_c26_c_fa2));
    FA fa_111(.A(stage0_r9_c17), .B(stage0_r10_c16), .C(stage0_r11_c15), .So(stage1_c26_s_fa3), .Co(stage1_c26_c_fa3));
    FA fa_112(.A(stage0_r12_c14), .B(stage0_r13_c13), .C(stage0_r14_c12), .So(stage1_c26_s_fa4), .Co(stage1_c26_c_fa4));
    FA fa_113(.A(stage0_r15_c11), .B(stage0_r16_c10), .C(stage0_r17_c9), .So(stage1_c26_s_fa5), .Co(stage1_c26_c_fa5));
    FA fa_114(.A(stage0_r18_c8), .B(stage0_r19_c7), .C(stage0_r20_c6), .So(stage1_c26_s_fa6), .Co(stage1_c26_c_fa6));
    FA fa_115(.A(stage0_r21_c5), .B(stage0_r22_c4), .C(stage0_r23_c3), .So(stage1_c26_s_fa7), .Co(stage1_c26_c_fa7));
    FA fa_116(.A(stage0_r24_c2), .B(stage0_r25_c1), .C(stage0_r26_c0), .So(stage1_c26_s_fa8), .Co(stage1_c26_c_fa8));
    FA fa_117(.A(stage0_r0_c27), .B(stage0_r1_c26), .C(stage0_r2_c25), .So(stage1_c27_s_fa0), .Co(stage1_c27_c_fa0));
    FA fa_118(.A(stage0_r3_c24), .B(stage0_r4_c23), .C(stage0_r5_c22), .So(stage1_c27_s_fa1), .Co(stage1_c27_c_fa1));
    FA fa_119(.A(stage0_r6_c21), .B(stage0_r7_c20), .C(stage0_r8_c19), .So(stage1_c27_s_fa2), .Co(stage1_c27_c_fa2));
    FA fa_120(.A(stage0_r9_c18), .B(stage0_r10_c17), .C(stage0_r11_c16), .So(stage1_c27_s_fa3), .Co(stage1_c27_c_fa3));
    FA fa_121(.A(stage0_r12_c15), .B(stage0_r13_c14), .C(stage0_r14_c13), .So(stage1_c27_s_fa4), .Co(stage1_c27_c_fa4));
    FA fa_122(.A(stage0_r15_c12), .B(stage0_r16_c11), .C(stage0_r17_c10), .So(stage1_c27_s_fa5), .Co(stage1_c27_c_fa5));
    FA fa_123(.A(stage0_r18_c9), .B(stage0_r19_c8), .C(stage0_r20_c7), .So(stage1_c27_s_fa6), .Co(stage1_c27_c_fa6));
    FA fa_124(.A(stage0_r21_c6), .B(stage0_r22_c5), .C(stage0_r23_c4), .So(stage1_c27_s_fa7), .Co(stage1_c27_c_fa7));
    FA fa_125(.A(stage0_r24_c3), .B(stage0_r25_c2), .C(stage0_r26_c1), .So(stage1_c27_s_fa8), .Co(stage1_c27_c_fa8));
    FA fa_126(.A(stage0_r0_c28), .B(stage0_r1_c27), .C(stage0_r2_c26), .So(stage1_c28_s_fa0), .Co(stage1_c28_c_fa0));
    FA fa_127(.A(stage0_r3_c25), .B(stage0_r4_c24), .C(stage0_r5_c23), .So(stage1_c28_s_fa1), .Co(stage1_c28_c_fa1));
    FA fa_128(.A(stage0_r6_c22), .B(stage0_r7_c21), .C(stage0_r8_c20), .So(stage1_c28_s_fa2), .Co(stage1_c28_c_fa2));
    FA fa_129(.A(stage0_r9_c19), .B(stage0_r10_c18), .C(stage0_r11_c17), .So(stage1_c28_s_fa3), .Co(stage1_c28_c_fa3));
    FA fa_130(.A(stage0_r12_c16), .B(stage0_r13_c15), .C(stage0_r14_c14), .So(stage1_c28_s_fa4), .Co(stage1_c28_c_fa4));
    FA fa_131(.A(stage0_r15_c13), .B(stage0_r16_c12), .C(stage0_r17_c11), .So(stage1_c28_s_fa5), .Co(stage1_c28_c_fa5));
    FA fa_132(.A(stage0_r18_c10), .B(stage0_r19_c9), .C(stage0_r20_c8), .So(stage1_c28_s_fa6), .Co(stage1_c28_c_fa6));
    FA fa_133(.A(stage0_r21_c7), .B(stage0_r22_c6), .C(stage0_r23_c5), .So(stage1_c28_s_fa7), .Co(stage1_c28_c_fa7));
    FA fa_134(.A(stage0_r24_c4), .B(stage0_r25_c3), .C(stage0_r26_c2), .So(stage1_c28_s_fa8), .Co(stage1_c28_c_fa8));
    HA ha_9(.A(stage0_r27_c1), .B(stage0_r28_c0), .So(stage1_c28_s_ha0), .Co(stage1_c28_c_ha0));
    FA fa_135(.A(stage0_r0_c29), .B(stage0_r1_c28), .C(stage0_r2_c27), .So(stage1_c29_s_fa0), .Co(stage1_c29_c_fa0));
    FA fa_136(.A(stage0_r3_c26), .B(stage0_r4_c25), .C(stage0_r5_c24), .So(stage1_c29_s_fa1), .Co(stage1_c29_c_fa1));
    FA fa_137(.A(stage0_r6_c23), .B(stage0_r7_c22), .C(stage0_r8_c21), .So(stage1_c29_s_fa2), .Co(stage1_c29_c_fa2));
    FA fa_138(.A(stage0_r9_c20), .B(stage0_r10_c19), .C(stage0_r11_c18), .So(stage1_c29_s_fa3), .Co(stage1_c29_c_fa3));
    FA fa_139(.A(stage0_r12_c17), .B(stage0_r13_c16), .C(stage0_r14_c15), .So(stage1_c29_s_fa4), .Co(stage1_c29_c_fa4));
    FA fa_140(.A(stage0_r15_c14), .B(stage0_r16_c13), .C(stage0_r17_c12), .So(stage1_c29_s_fa5), .Co(stage1_c29_c_fa5));
    FA fa_141(.A(stage0_r18_c11), .B(stage0_r19_c10), .C(stage0_r20_c9), .So(stage1_c29_s_fa6), .Co(stage1_c29_c_fa6));
    FA fa_142(.A(stage0_r21_c8), .B(stage0_r22_c7), .C(stage0_r23_c6), .So(stage1_c29_s_fa7), .Co(stage1_c29_c_fa7));
    FA fa_143(.A(stage0_r24_c5), .B(stage0_r25_c4), .C(stage0_r26_c3), .So(stage1_c29_s_fa8), .Co(stage1_c29_c_fa8));
    FA fa_144(.A(stage0_r27_c2), .B(stage0_r28_c1), .C(stage0_r29_c0), .So(stage1_c29_s_fa9), .Co(stage1_c29_c_fa9));
    FA fa_145(.A(stage0_r0_c30), .B(stage0_r1_c29), .C(stage0_r2_c28), .So(stage1_c30_s_fa0), .Co(stage1_c30_c_fa0));
    FA fa_146(.A(stage0_r3_c27), .B(stage0_r4_c26), .C(stage0_r5_c25), .So(stage1_c30_s_fa1), .Co(stage1_c30_c_fa1));
    FA fa_147(.A(stage0_r6_c24), .B(stage0_r7_c23), .C(stage0_r8_c22), .So(stage1_c30_s_fa2), .Co(stage1_c30_c_fa2));
    FA fa_148(.A(stage0_r9_c21), .B(stage0_r10_c20), .C(stage0_r11_c19), .So(stage1_c30_s_fa3), .Co(stage1_c30_c_fa3));
    FA fa_149(.A(stage0_r12_c18), .B(stage0_r13_c17), .C(stage0_r14_c16), .So(stage1_c30_s_fa4), .Co(stage1_c30_c_fa4));
    FA fa_150(.A(stage0_r15_c15), .B(stage0_r16_c14), .C(stage0_r17_c13), .So(stage1_c30_s_fa5), .Co(stage1_c30_c_fa5));
    FA fa_151(.A(stage0_r18_c12), .B(stage0_r19_c11), .C(stage0_r20_c10), .So(stage1_c30_s_fa6), .Co(stage1_c30_c_fa6));
    FA fa_152(.A(stage0_r21_c9), .B(stage0_r22_c8), .C(stage0_r23_c7), .So(stage1_c30_s_fa7), .Co(stage1_c30_c_fa7));
    FA fa_153(.A(stage0_r24_c6), .B(stage0_r25_c5), .C(stage0_r26_c4), .So(stage1_c30_s_fa8), .Co(stage1_c30_c_fa8));
    FA fa_154(.A(stage0_r27_c3), .B(stage0_r28_c2), .C(stage0_r29_c1), .So(stage1_c30_s_fa9), .Co(stage1_c30_c_fa9));
    FA fa_155(.A(stage0_r0_c31), .B(stage0_r1_c30), .C(stage0_r2_c29), .So(stage1_c31_s_fa0), .Co(stage1_c31_c_fa0));
    FA fa_156(.A(stage0_r3_c28), .B(stage0_r4_c27), .C(stage0_r5_c26), .So(stage1_c31_s_fa1), .Co(stage1_c31_c_fa1));
    FA fa_157(.A(stage0_r6_c25), .B(stage0_r7_c24), .C(stage0_r8_c23), .So(stage1_c31_s_fa2), .Co(stage1_c31_c_fa2));
    FA fa_158(.A(stage0_r9_c22), .B(stage0_r10_c21), .C(stage0_r11_c20), .So(stage1_c31_s_fa3), .Co(stage1_c31_c_fa3));
    FA fa_159(.A(stage0_r12_c19), .B(stage0_r13_c18), .C(stage0_r14_c17), .So(stage1_c31_s_fa4), .Co(stage1_c31_c_fa4));
    FA fa_160(.A(stage0_r15_c16), .B(stage0_r16_c15), .C(stage0_r17_c14), .So(stage1_c31_s_fa5), .Co(stage1_c31_c_fa5));
    FA fa_161(.A(stage0_r18_c13), .B(stage0_r19_c12), .C(stage0_r20_c11), .So(stage1_c31_s_fa6), .Co(stage1_c31_c_fa6));
    FA fa_162(.A(stage0_r21_c10), .B(stage0_r22_c9), .C(stage0_r23_c8), .So(stage1_c31_s_fa7), .Co(stage1_c31_c_fa7));
    FA fa_163(.A(stage0_r24_c7), .B(stage0_r25_c6), .C(stage0_r26_c5), .So(stage1_c31_s_fa8), .Co(stage1_c31_c_fa8));
    FA fa_164(.A(stage0_r27_c4), .B(stage0_r28_c3), .C(stage0_r29_c2), .So(stage1_c31_s_fa9), .Co(stage1_c31_c_fa9));
    HA ha_10(.A(stage0_r30_c1), .B(stage0_r31_c0), .So(stage1_c31_s_ha0), .Co(stage1_c31_c_ha0));
    FA fa_165(.A(stage0_r0_c32), .B(stage0_r1_c31), .C(stage0_r2_c30), .So(stage1_c32_s_fa0), .Co(stage1_c32_c_fa0));
    FA fa_166(.A(stage0_r3_c29), .B(stage0_r4_c28), .C(stage0_r5_c27), .So(stage1_c32_s_fa1), .Co(stage1_c32_c_fa1));
    FA fa_167(.A(stage0_r6_c26), .B(stage0_r7_c25), .C(stage0_r8_c24), .So(stage1_c32_s_fa2), .Co(stage1_c32_c_fa2));
    FA fa_168(.A(stage0_r9_c23), .B(stage0_r10_c22), .C(stage0_r11_c21), .So(stage1_c32_s_fa3), .Co(stage1_c32_c_fa3));
    FA fa_169(.A(stage0_r12_c20), .B(stage0_r13_c19), .C(stage0_r14_c18), .So(stage1_c32_s_fa4), .Co(stage1_c32_c_fa4));
    FA fa_170(.A(stage0_r15_c17), .B(stage0_r16_c16), .C(stage0_r17_c15), .So(stage1_c32_s_fa5), .Co(stage1_c32_c_fa5));
    FA fa_171(.A(stage0_r18_c14), .B(stage0_r19_c13), .C(stage0_r20_c12), .So(stage1_c32_s_fa6), .Co(stage1_c32_c_fa6));
    FA fa_172(.A(stage0_r21_c11), .B(stage0_r22_c10), .C(stage0_r23_c9), .So(stage1_c32_s_fa7), .Co(stage1_c32_c_fa7));
    FA fa_173(.A(stage0_r24_c8), .B(stage0_r25_c7), .C(stage0_r26_c6), .So(stage1_c32_s_fa8), .Co(stage1_c32_c_fa8));
    FA fa_174(.A(stage0_r27_c5), .B(stage0_r28_c4), .C(stage0_r29_c3), .So(stage1_c32_s_fa9), .Co(stage1_c32_c_fa9));
    FA fa_175(.A(stage0_r30_c2), .B(stage0_r31_c1), .C(stage0_r32_c0), .So(stage1_c32_s_fa10), .Co(stage1_c32_c_fa10));
    FA fa_176(.A(stage0_r0_c33), .B(stage0_r1_c32), .C(stage0_r2_c31), .So(stage1_c33_s_fa0), .Co(stage1_c33_c_fa0));
    FA fa_177(.A(stage0_r3_c30), .B(stage0_r4_c29), .C(stage0_r5_c28), .So(stage1_c33_s_fa1), .Co(stage1_c33_c_fa1));
    FA fa_178(.A(stage0_r6_c27), .B(stage0_r7_c26), .C(stage0_r8_c25), .So(stage1_c33_s_fa2), .Co(stage1_c33_c_fa2));
    FA fa_179(.A(stage0_r9_c24), .B(stage0_r10_c23), .C(stage0_r11_c22), .So(stage1_c33_s_fa3), .Co(stage1_c33_c_fa3));
    FA fa_180(.A(stage0_r12_c21), .B(stage0_r13_c20), .C(stage0_r14_c19), .So(stage1_c33_s_fa4), .Co(stage1_c33_c_fa4));
    FA fa_181(.A(stage0_r15_c18), .B(stage0_r16_c17), .C(stage0_r17_c16), .So(stage1_c33_s_fa5), .Co(stage1_c33_c_fa5));
    FA fa_182(.A(stage0_r18_c15), .B(stage0_r19_c14), .C(stage0_r20_c13), .So(stage1_c33_s_fa6), .Co(stage1_c33_c_fa6));
    FA fa_183(.A(stage0_r21_c12), .B(stage0_r22_c11), .C(stage0_r23_c10), .So(stage1_c33_s_fa7), .Co(stage1_c33_c_fa7));
    FA fa_184(.A(stage0_r24_c9), .B(stage0_r25_c8), .C(stage0_r26_c7), .So(stage1_c33_s_fa8), .Co(stage1_c33_c_fa8));
    FA fa_185(.A(stage0_r27_c6), .B(stage0_r28_c5), .C(stage0_r29_c4), .So(stage1_c33_s_fa9), .Co(stage1_c33_c_fa9));
    FA fa_186(.A(stage0_r30_c3), .B(stage0_r31_c2), .C(stage0_r32_c1), .So(stage1_c33_s_fa10), .Co(stage1_c33_c_fa10));
    FA fa_187(.A(stage0_r0_c34), .B(stage0_r1_c33), .C(stage0_r2_c32), .So(stage1_c34_s_fa0), .Co(stage1_c34_c_fa0));
    FA fa_188(.A(stage0_r3_c31), .B(stage0_r4_c30), .C(stage0_r5_c29), .So(stage1_c34_s_fa1), .Co(stage1_c34_c_fa1));
    FA fa_189(.A(stage0_r6_c28), .B(stage0_r7_c27), .C(stage0_r8_c26), .So(stage1_c34_s_fa2), .Co(stage1_c34_c_fa2));
    FA fa_190(.A(stage0_r9_c25), .B(stage0_r10_c24), .C(stage0_r11_c23), .So(stage1_c34_s_fa3), .Co(stage1_c34_c_fa3));
    FA fa_191(.A(stage0_r12_c22), .B(stage0_r13_c21), .C(stage0_r14_c20), .So(stage1_c34_s_fa4), .Co(stage1_c34_c_fa4));
    FA fa_192(.A(stage0_r15_c19), .B(stage0_r16_c18), .C(stage0_r17_c17), .So(stage1_c34_s_fa5), .Co(stage1_c34_c_fa5));
    FA fa_193(.A(stage0_r18_c16), .B(stage0_r19_c15), .C(stage0_r20_c14), .So(stage1_c34_s_fa6), .Co(stage1_c34_c_fa6));
    FA fa_194(.A(stage0_r21_c13), .B(stage0_r22_c12), .C(stage0_r23_c11), .So(stage1_c34_s_fa7), .Co(stage1_c34_c_fa7));
    FA fa_195(.A(stage0_r24_c10), .B(stage0_r25_c9), .C(stage0_r26_c8), .So(stage1_c34_s_fa8), .Co(stage1_c34_c_fa8));
    FA fa_196(.A(stage0_r27_c7), .B(stage0_r28_c6), .C(stage0_r29_c5), .So(stage1_c34_s_fa9), .Co(stage1_c34_c_fa9));
    FA fa_197(.A(stage0_r30_c4), .B(stage0_r31_c3), .C(stage0_r32_c2), .So(stage1_c34_s_fa10), .Co(stage1_c34_c_fa10));
    HA ha_11(.A(stage0_r33_c1), .B(stage0_r34_c0), .So(stage1_c34_s_ha0), .Co(stage1_c34_c_ha0));
    FA fa_198(.A(stage0_r0_c35), .B(stage0_r1_c34), .C(stage0_r2_c33), .So(stage1_c35_s_fa0), .Co(stage1_c35_c_fa0));
    FA fa_199(.A(stage0_r3_c32), .B(stage0_r4_c31), .C(stage0_r5_c30), .So(stage1_c35_s_fa1), .Co(stage1_c35_c_fa1));
    FA fa_200(.A(stage0_r6_c29), .B(stage0_r7_c28), .C(stage0_r8_c27), .So(stage1_c35_s_fa2), .Co(stage1_c35_c_fa2));
    FA fa_201(.A(stage0_r9_c26), .B(stage0_r10_c25), .C(stage0_r11_c24), .So(stage1_c35_s_fa3), .Co(stage1_c35_c_fa3));
    FA fa_202(.A(stage0_r12_c23), .B(stage0_r13_c22), .C(stage0_r14_c21), .So(stage1_c35_s_fa4), .Co(stage1_c35_c_fa4));
    FA fa_203(.A(stage0_r15_c20), .B(stage0_r16_c19), .C(stage0_r17_c18), .So(stage1_c35_s_fa5), .Co(stage1_c35_c_fa5));
    FA fa_204(.A(stage0_r18_c17), .B(stage0_r19_c16), .C(stage0_r20_c15), .So(stage1_c35_s_fa6), .Co(stage1_c35_c_fa6));
    FA fa_205(.A(stage0_r21_c14), .B(stage0_r22_c13), .C(stage0_r23_c12), .So(stage1_c35_s_fa7), .Co(stage1_c35_c_fa7));
    FA fa_206(.A(stage0_r24_c11), .B(stage0_r25_c10), .C(stage0_r26_c9), .So(stage1_c35_s_fa8), .Co(stage1_c35_c_fa8));
    FA fa_207(.A(stage0_r27_c8), .B(stage0_r28_c7), .C(stage0_r29_c6), .So(stage1_c35_s_fa9), .Co(stage1_c35_c_fa9));
    FA fa_208(.A(stage0_r30_c5), .B(stage0_r31_c4), .C(stage0_r32_c3), .So(stage1_c35_s_fa10), .Co(stage1_c35_c_fa10));
    FA fa_209(.A(stage0_r33_c2), .B(stage0_r34_c1), .C(stage0_r35_c0), .So(stage1_c35_s_fa11), .Co(stage1_c35_c_fa11));
    FA fa_210(.A(stage0_r0_c36), .B(stage0_r1_c35), .C(stage0_r2_c34), .So(stage1_c36_s_fa0), .Co(stage1_c36_c_fa0));
    FA fa_211(.A(stage0_r3_c33), .B(stage0_r4_c32), .C(stage0_r5_c31), .So(stage1_c36_s_fa1), .Co(stage1_c36_c_fa1));
    FA fa_212(.A(stage0_r6_c30), .B(stage0_r7_c29), .C(stage0_r8_c28), .So(stage1_c36_s_fa2), .Co(stage1_c36_c_fa2));
    FA fa_213(.A(stage0_r9_c27), .B(stage0_r10_c26), .C(stage0_r11_c25), .So(stage1_c36_s_fa3), .Co(stage1_c36_c_fa3));
    FA fa_214(.A(stage0_r12_c24), .B(stage0_r13_c23), .C(stage0_r14_c22), .So(stage1_c36_s_fa4), .Co(stage1_c36_c_fa4));
    FA fa_215(.A(stage0_r15_c21), .B(stage0_r16_c20), .C(stage0_r17_c19), .So(stage1_c36_s_fa5), .Co(stage1_c36_c_fa5));
    FA fa_216(.A(stage0_r18_c18), .B(stage0_r19_c17), .C(stage0_r20_c16), .So(stage1_c36_s_fa6), .Co(stage1_c36_c_fa6));
    FA fa_217(.A(stage0_r21_c15), .B(stage0_r22_c14), .C(stage0_r23_c13), .So(stage1_c36_s_fa7), .Co(stage1_c36_c_fa7));
    FA fa_218(.A(stage0_r24_c12), .B(stage0_r25_c11), .C(stage0_r26_c10), .So(stage1_c36_s_fa8), .Co(stage1_c36_c_fa8));
    FA fa_219(.A(stage0_r27_c9), .B(stage0_r28_c8), .C(stage0_r29_c7), .So(stage1_c36_s_fa9), .Co(stage1_c36_c_fa9));
    FA fa_220(.A(stage0_r30_c6), .B(stage0_r31_c5), .C(stage0_r32_c4), .So(stage1_c36_s_fa10), .Co(stage1_c36_c_fa10));
    FA fa_221(.A(stage0_r33_c3), .B(stage0_r34_c2), .C(stage0_r35_c1), .So(stage1_c36_s_fa11), .Co(stage1_c36_c_fa11));
    FA fa_222(.A(stage0_r0_c37), .B(stage0_r1_c36), .C(stage0_r2_c35), .So(stage1_c37_s_fa0), .Co(stage1_c37_c_fa0));
    FA fa_223(.A(stage0_r3_c34), .B(stage0_r4_c33), .C(stage0_r5_c32), .So(stage1_c37_s_fa1), .Co(stage1_c37_c_fa1));
    FA fa_224(.A(stage0_r6_c31), .B(stage0_r7_c30), .C(stage0_r8_c29), .So(stage1_c37_s_fa2), .Co(stage1_c37_c_fa2));
    FA fa_225(.A(stage0_r9_c28), .B(stage0_r10_c27), .C(stage0_r11_c26), .So(stage1_c37_s_fa3), .Co(stage1_c37_c_fa3));
    FA fa_226(.A(stage0_r12_c25), .B(stage0_r13_c24), .C(stage0_r14_c23), .So(stage1_c37_s_fa4), .Co(stage1_c37_c_fa4));
    FA fa_227(.A(stage0_r15_c22), .B(stage0_r16_c21), .C(stage0_r17_c20), .So(stage1_c37_s_fa5), .Co(stage1_c37_c_fa5));
    FA fa_228(.A(stage0_r18_c19), .B(stage0_r19_c18), .C(stage0_r20_c17), .So(stage1_c37_s_fa6), .Co(stage1_c37_c_fa6));
    FA fa_229(.A(stage0_r21_c16), .B(stage0_r22_c15), .C(stage0_r23_c14), .So(stage1_c37_s_fa7), .Co(stage1_c37_c_fa7));
    FA fa_230(.A(stage0_r24_c13), .B(stage0_r25_c12), .C(stage0_r26_c11), .So(stage1_c37_s_fa8), .Co(stage1_c37_c_fa8));
    FA fa_231(.A(stage0_r27_c10), .B(stage0_r28_c9), .C(stage0_r29_c8), .So(stage1_c37_s_fa9), .Co(stage1_c37_c_fa9));
    FA fa_232(.A(stage0_r30_c7), .B(stage0_r31_c6), .C(stage0_r32_c5), .So(stage1_c37_s_fa10), .Co(stage1_c37_c_fa10));
    FA fa_233(.A(stage0_r33_c4), .B(stage0_r34_c3), .C(stage0_r35_c2), .So(stage1_c37_s_fa11), .Co(stage1_c37_c_fa11));
    HA ha_12(.A(stage0_r36_c1), .B(stage0_r37_c0), .So(stage1_c37_s_ha0), .Co(stage1_c37_c_ha0));
    FA fa_234(.A(stage0_r0_c38), .B(stage0_r1_c37), .C(stage0_r2_c36), .So(stage1_c38_s_fa0), .Co(stage1_c38_c_fa0));
    FA fa_235(.A(stage0_r3_c35), .B(stage0_r4_c34), .C(stage0_r5_c33), .So(stage1_c38_s_fa1), .Co(stage1_c38_c_fa1));
    FA fa_236(.A(stage0_r6_c32), .B(stage0_r7_c31), .C(stage0_r8_c30), .So(stage1_c38_s_fa2), .Co(stage1_c38_c_fa2));
    FA fa_237(.A(stage0_r9_c29), .B(stage0_r10_c28), .C(stage0_r11_c27), .So(stage1_c38_s_fa3), .Co(stage1_c38_c_fa3));
    FA fa_238(.A(stage0_r12_c26), .B(stage0_r13_c25), .C(stage0_r14_c24), .So(stage1_c38_s_fa4), .Co(stage1_c38_c_fa4));
    FA fa_239(.A(stage0_r15_c23), .B(stage0_r16_c22), .C(stage0_r17_c21), .So(stage1_c38_s_fa5), .Co(stage1_c38_c_fa5));
    FA fa_240(.A(stage0_r18_c20), .B(stage0_r19_c19), .C(stage0_r20_c18), .So(stage1_c38_s_fa6), .Co(stage1_c38_c_fa6));
    FA fa_241(.A(stage0_r21_c17), .B(stage0_r22_c16), .C(stage0_r23_c15), .So(stage1_c38_s_fa7), .Co(stage1_c38_c_fa7));
    FA fa_242(.A(stage0_r24_c14), .B(stage0_r25_c13), .C(stage0_r26_c12), .So(stage1_c38_s_fa8), .Co(stage1_c38_c_fa8));
    FA fa_243(.A(stage0_r27_c11), .B(stage0_r28_c10), .C(stage0_r29_c9), .So(stage1_c38_s_fa9), .Co(stage1_c38_c_fa9));
    FA fa_244(.A(stage0_r30_c8), .B(stage0_r31_c7), .C(stage0_r32_c6), .So(stage1_c38_s_fa10), .Co(stage1_c38_c_fa10));
    FA fa_245(.A(stage0_r33_c5), .B(stage0_r34_c4), .C(stage0_r35_c3), .So(stage1_c38_s_fa11), .Co(stage1_c38_c_fa11));
    FA fa_246(.A(stage0_r36_c2), .B(stage0_r37_c1), .C(stage0_r38_c0), .So(stage1_c38_s_fa12), .Co(stage1_c38_c_fa12));
    FA fa_247(.A(stage0_r0_c39), .B(stage0_r1_c38), .C(stage0_r2_c37), .So(stage1_c39_s_fa0), .Co(stage1_c39_c_fa0));
    FA fa_248(.A(stage0_r3_c36), .B(stage0_r4_c35), .C(stage0_r5_c34), .So(stage1_c39_s_fa1), .Co(stage1_c39_c_fa1));
    FA fa_249(.A(stage0_r6_c33), .B(stage0_r7_c32), .C(stage0_r8_c31), .So(stage1_c39_s_fa2), .Co(stage1_c39_c_fa2));
    FA fa_250(.A(stage0_r9_c30), .B(stage0_r10_c29), .C(stage0_r11_c28), .So(stage1_c39_s_fa3), .Co(stage1_c39_c_fa3));
    FA fa_251(.A(stage0_r12_c27), .B(stage0_r13_c26), .C(stage0_r14_c25), .So(stage1_c39_s_fa4), .Co(stage1_c39_c_fa4));
    FA fa_252(.A(stage0_r15_c24), .B(stage0_r16_c23), .C(stage0_r17_c22), .So(stage1_c39_s_fa5), .Co(stage1_c39_c_fa5));
    FA fa_253(.A(stage0_r18_c21), .B(stage0_r19_c20), .C(stage0_r20_c19), .So(stage1_c39_s_fa6), .Co(stage1_c39_c_fa6));
    FA fa_254(.A(stage0_r21_c18), .B(stage0_r22_c17), .C(stage0_r23_c16), .So(stage1_c39_s_fa7), .Co(stage1_c39_c_fa7));
    FA fa_255(.A(stage0_r24_c15), .B(stage0_r25_c14), .C(stage0_r26_c13), .So(stage1_c39_s_fa8), .Co(stage1_c39_c_fa8));
    FA fa_256(.A(stage0_r27_c12), .B(stage0_r28_c11), .C(stage0_r29_c10), .So(stage1_c39_s_fa9), .Co(stage1_c39_c_fa9));
    FA fa_257(.A(stage0_r30_c9), .B(stage0_r31_c8), .C(stage0_r32_c7), .So(stage1_c39_s_fa10), .Co(stage1_c39_c_fa10));
    FA fa_258(.A(stage0_r33_c6), .B(stage0_r34_c5), .C(stage0_r35_c4), .So(stage1_c39_s_fa11), .Co(stage1_c39_c_fa11));
    FA fa_259(.A(stage0_r36_c3), .B(stage0_r37_c2), .C(stage0_r38_c1), .So(stage1_c39_s_fa12), .Co(stage1_c39_c_fa12));
    FA fa_260(.A(stage0_r0_c40), .B(stage0_r1_c39), .C(stage0_r2_c38), .So(stage1_c40_s_fa0), .Co(stage1_c40_c_fa0));
    FA fa_261(.A(stage0_r3_c37), .B(stage0_r4_c36), .C(stage0_r5_c35), .So(stage1_c40_s_fa1), .Co(stage1_c40_c_fa1));
    FA fa_262(.A(stage0_r6_c34), .B(stage0_r7_c33), .C(stage0_r8_c32), .So(stage1_c40_s_fa2), .Co(stage1_c40_c_fa2));
    FA fa_263(.A(stage0_r9_c31), .B(stage0_r10_c30), .C(stage0_r11_c29), .So(stage1_c40_s_fa3), .Co(stage1_c40_c_fa3));
    FA fa_264(.A(stage0_r12_c28), .B(stage0_r13_c27), .C(stage0_r14_c26), .So(stage1_c40_s_fa4), .Co(stage1_c40_c_fa4));
    FA fa_265(.A(stage0_r15_c25), .B(stage0_r16_c24), .C(stage0_r17_c23), .So(stage1_c40_s_fa5), .Co(stage1_c40_c_fa5));
    FA fa_266(.A(stage0_r18_c22), .B(stage0_r19_c21), .C(stage0_r20_c20), .So(stage1_c40_s_fa6), .Co(stage1_c40_c_fa6));
    FA fa_267(.A(stage0_r21_c19), .B(stage0_r22_c18), .C(stage0_r23_c17), .So(stage1_c40_s_fa7), .Co(stage1_c40_c_fa7));
    FA fa_268(.A(stage0_r24_c16), .B(stage0_r25_c15), .C(stage0_r26_c14), .So(stage1_c40_s_fa8), .Co(stage1_c40_c_fa8));
    FA fa_269(.A(stage0_r27_c13), .B(stage0_r28_c12), .C(stage0_r29_c11), .So(stage1_c40_s_fa9), .Co(stage1_c40_c_fa9));
    FA fa_270(.A(stage0_r30_c10), .B(stage0_r31_c9), .C(stage0_r32_c8), .So(stage1_c40_s_fa10), .Co(stage1_c40_c_fa10));
    FA fa_271(.A(stage0_r33_c7), .B(stage0_r34_c6), .C(stage0_r35_c5), .So(stage1_c40_s_fa11), .Co(stage1_c40_c_fa11));
    FA fa_272(.A(stage0_r36_c4), .B(stage0_r37_c3), .C(stage0_r38_c2), .So(stage1_c40_s_fa12), .Co(stage1_c40_c_fa12));
    HA ha_13(.A(stage0_r39_c1), .B(stage0_r40_c0), .So(stage1_c40_s_ha0), .Co(stage1_c40_c_ha0));
    FA fa_273(.A(stage0_r1_c40), .B(stage0_r2_c39), .C(stage0_r3_c38), .So(stage1_c41_s_fa0), .Co(stage1_c41_c_fa0));
    FA fa_274(.A(stage0_r4_c37), .B(stage0_r5_c36), .C(stage0_r6_c35), .So(stage1_c41_s_fa1), .Co(stage1_c41_c_fa1));
    FA fa_275(.A(stage0_r7_c34), .B(stage0_r8_c33), .C(stage0_r9_c32), .So(stage1_c41_s_fa2), .Co(stage1_c41_c_fa2));
    FA fa_276(.A(stage0_r10_c31), .B(stage0_r11_c30), .C(stage0_r12_c29), .So(stage1_c41_s_fa3), .Co(stage1_c41_c_fa3));
    FA fa_277(.A(stage0_r13_c28), .B(stage0_r14_c27), .C(stage0_r15_c26), .So(stage1_c41_s_fa4), .Co(stage1_c41_c_fa4));
    FA fa_278(.A(stage0_r16_c25), .B(stage0_r17_c24), .C(stage0_r18_c23), .So(stage1_c41_s_fa5), .Co(stage1_c41_c_fa5));
    FA fa_279(.A(stage0_r19_c22), .B(stage0_r20_c21), .C(stage0_r21_c20), .So(stage1_c41_s_fa6), .Co(stage1_c41_c_fa6));
    FA fa_280(.A(stage0_r22_c19), .B(stage0_r23_c18), .C(stage0_r24_c17), .So(stage1_c41_s_fa7), .Co(stage1_c41_c_fa7));
    FA fa_281(.A(stage0_r25_c16), .B(stage0_r26_c15), .C(stage0_r27_c14), .So(stage1_c41_s_fa8), .Co(stage1_c41_c_fa8));
    FA fa_282(.A(stage0_r28_c13), .B(stage0_r29_c12), .C(stage0_r30_c11), .So(stage1_c41_s_fa9), .Co(stage1_c41_c_fa9));
    FA fa_283(.A(stage0_r31_c10), .B(stage0_r32_c9), .C(stage0_r33_c8), .So(stage1_c41_s_fa10), .Co(stage1_c41_c_fa10));
    FA fa_284(.A(stage0_r34_c7), .B(stage0_r35_c6), .C(stage0_r36_c5), .So(stage1_c41_s_fa11), .Co(stage1_c41_c_fa11));
    FA fa_285(.A(stage0_r37_c4), .B(stage0_r38_c3), .C(stage0_r39_c2), .So(stage1_c41_s_fa12), .Co(stage1_c41_c_fa12));
    HA ha_14(.A(stage0_r40_c1), .B(stage0_r41_c0), .So(stage1_c41_s_ha0), .Co(stage1_c41_c_ha0));
    FA fa_286(.A(stage0_r2_c40), .B(stage0_r3_c39), .C(stage0_r4_c38), .So(stage1_c42_s_fa0), .Co(stage1_c42_c_fa0));
    FA fa_287(.A(stage0_r5_c37), .B(stage0_r6_c36), .C(stage0_r7_c35), .So(stage1_c42_s_fa1), .Co(stage1_c42_c_fa1));
    FA fa_288(.A(stage0_r8_c34), .B(stage0_r9_c33), .C(stage0_r10_c32), .So(stage1_c42_s_fa2), .Co(stage1_c42_c_fa2));
    FA fa_289(.A(stage0_r11_c31), .B(stage0_r12_c30), .C(stage0_r13_c29), .So(stage1_c42_s_fa3), .Co(stage1_c42_c_fa3));
    FA fa_290(.A(stage0_r14_c28), .B(stage0_r15_c27), .C(stage0_r16_c26), .So(stage1_c42_s_fa4), .Co(stage1_c42_c_fa4));
    FA fa_291(.A(stage0_r17_c25), .B(stage0_r18_c24), .C(stage0_r19_c23), .So(stage1_c42_s_fa5), .Co(stage1_c42_c_fa5));
    FA fa_292(.A(stage0_r20_c22), .B(stage0_r21_c21), .C(stage0_r22_c20), .So(stage1_c42_s_fa6), .Co(stage1_c42_c_fa6));
    FA fa_293(.A(stage0_r23_c19), .B(stage0_r24_c18), .C(stage0_r25_c17), .So(stage1_c42_s_fa7), .Co(stage1_c42_c_fa7));
    FA fa_294(.A(stage0_r26_c16), .B(stage0_r27_c15), .C(stage0_r28_c14), .So(stage1_c42_s_fa8), .Co(stage1_c42_c_fa8));
    FA fa_295(.A(stage0_r29_c13), .B(stage0_r30_c12), .C(stage0_r31_c11), .So(stage1_c42_s_fa9), .Co(stage1_c42_c_fa9));
    FA fa_296(.A(stage0_r32_c10), .B(stage0_r33_c9), .C(stage0_r34_c8), .So(stage1_c42_s_fa10), .Co(stage1_c42_c_fa10));
    FA fa_297(.A(stage0_r35_c7), .B(stage0_r36_c6), .C(stage0_r37_c5), .So(stage1_c42_s_fa11), .Co(stage1_c42_c_fa11));
    FA fa_298(.A(stage0_r38_c4), .B(stage0_r39_c3), .C(stage0_r40_c2), .So(stage1_c42_s_fa12), .Co(stage1_c42_c_fa12));
    HA ha_15(.A(stage0_r41_c1), .B(stage0_r42_c0), .So(stage1_c42_s_ha0), .Co(stage1_c42_c_ha0));
    FA fa_299(.A(stage0_r3_c40), .B(stage0_r4_c39), .C(stage0_r5_c38), .So(stage1_c43_s_fa0), .Co(stage1_c43_c_fa0));
    FA fa_300(.A(stage0_r6_c37), .B(stage0_r7_c36), .C(stage0_r8_c35), .So(stage1_c43_s_fa1), .Co(stage1_c43_c_fa1));
    FA fa_301(.A(stage0_r9_c34), .B(stage0_r10_c33), .C(stage0_r11_c32), .So(stage1_c43_s_fa2), .Co(stage1_c43_c_fa2));
    FA fa_302(.A(stage0_r12_c31), .B(stage0_r13_c30), .C(stage0_r14_c29), .So(stage1_c43_s_fa3), .Co(stage1_c43_c_fa3));
    FA fa_303(.A(stage0_r15_c28), .B(stage0_r16_c27), .C(stage0_r17_c26), .So(stage1_c43_s_fa4), .Co(stage1_c43_c_fa4));
    FA fa_304(.A(stage0_r18_c25), .B(stage0_r19_c24), .C(stage0_r20_c23), .So(stage1_c43_s_fa5), .Co(stage1_c43_c_fa5));
    FA fa_305(.A(stage0_r21_c22), .B(stage0_r22_c21), .C(stage0_r23_c20), .So(stage1_c43_s_fa6), .Co(stage1_c43_c_fa6));
    FA fa_306(.A(stage0_r24_c19), .B(stage0_r25_c18), .C(stage0_r26_c17), .So(stage1_c43_s_fa7), .Co(stage1_c43_c_fa7));
    FA fa_307(.A(stage0_r27_c16), .B(stage0_r28_c15), .C(stage0_r29_c14), .So(stage1_c43_s_fa8), .Co(stage1_c43_c_fa8));
    FA fa_308(.A(stage0_r30_c13), .B(stage0_r31_c12), .C(stage0_r32_c11), .So(stage1_c43_s_fa9), .Co(stage1_c43_c_fa9));
    FA fa_309(.A(stage0_r33_c10), .B(stage0_r34_c9), .C(stage0_r35_c8), .So(stage1_c43_s_fa10), .Co(stage1_c43_c_fa10));
    FA fa_310(.A(stage0_r36_c7), .B(stage0_r37_c6), .C(stage0_r38_c5), .So(stage1_c43_s_fa11), .Co(stage1_c43_c_fa11));
    FA fa_311(.A(stage0_r39_c4), .B(stage0_r40_c3), .C(stage0_r41_c2), .So(stage1_c43_s_fa12), .Co(stage1_c43_c_fa12));
    HA ha_16(.A(stage0_r42_c1), .B(stage0_r43_c0), .So(stage1_c43_s_ha0), .Co(stage1_c43_c_ha0));
    FA fa_312(.A(stage0_r4_c40), .B(stage0_r5_c39), .C(stage0_r6_c38), .So(stage1_c44_s_fa0), .Co(stage1_c44_c_fa0));
    FA fa_313(.A(stage0_r7_c37), .B(stage0_r8_c36), .C(stage0_r9_c35), .So(stage1_c44_s_fa1), .Co(stage1_c44_c_fa1));
    FA fa_314(.A(stage0_r10_c34), .B(stage0_r11_c33), .C(stage0_r12_c32), .So(stage1_c44_s_fa2), .Co(stage1_c44_c_fa2));
    FA fa_315(.A(stage0_r13_c31), .B(stage0_r14_c30), .C(stage0_r15_c29), .So(stage1_c44_s_fa3), .Co(stage1_c44_c_fa3));
    FA fa_316(.A(stage0_r16_c28), .B(stage0_r17_c27), .C(stage0_r18_c26), .So(stage1_c44_s_fa4), .Co(stage1_c44_c_fa4));
    FA fa_317(.A(stage0_r19_c25), .B(stage0_r20_c24), .C(stage0_r21_c23), .So(stage1_c44_s_fa5), .Co(stage1_c44_c_fa5));
    FA fa_318(.A(stage0_r22_c22), .B(stage0_r23_c21), .C(stage0_r24_c20), .So(stage1_c44_s_fa6), .Co(stage1_c44_c_fa6));
    FA fa_319(.A(stage0_r25_c19), .B(stage0_r26_c18), .C(stage0_r27_c17), .So(stage1_c44_s_fa7), .Co(stage1_c44_c_fa7));
    FA fa_320(.A(stage0_r28_c16), .B(stage0_r29_c15), .C(stage0_r30_c14), .So(stage1_c44_s_fa8), .Co(stage1_c44_c_fa8));
    FA fa_321(.A(stage0_r31_c13), .B(stage0_r32_c12), .C(stage0_r33_c11), .So(stage1_c44_s_fa9), .Co(stage1_c44_c_fa9));
    FA fa_322(.A(stage0_r34_c10), .B(stage0_r35_c9), .C(stage0_r36_c8), .So(stage1_c44_s_fa10), .Co(stage1_c44_c_fa10));
    FA fa_323(.A(stage0_r37_c7), .B(stage0_r38_c6), .C(stage0_r39_c5), .So(stage1_c44_s_fa11), .Co(stage1_c44_c_fa11));
    FA fa_324(.A(stage0_r40_c4), .B(stage0_r41_c3), .C(stage0_r42_c2), .So(stage1_c44_s_fa12), .Co(stage1_c44_c_fa12));
    HA ha_17(.A(stage0_r43_c1), .B(stage0_r44_c0), .So(stage1_c44_s_ha0), .Co(stage1_c44_c_ha0));
    FA fa_325(.A(stage0_r5_c40), .B(stage0_r6_c39), .C(stage0_r7_c38), .So(stage1_c45_s_fa0), .Co(stage1_c45_c_fa0));
    FA fa_326(.A(stage0_r8_c37), .B(stage0_r9_c36), .C(stage0_r10_c35), .So(stage1_c45_s_fa1), .Co(stage1_c45_c_fa1));
    FA fa_327(.A(stage0_r11_c34), .B(stage0_r12_c33), .C(stage0_r13_c32), .So(stage1_c45_s_fa2), .Co(stage1_c45_c_fa2));
    FA fa_328(.A(stage0_r14_c31), .B(stage0_r15_c30), .C(stage0_r16_c29), .So(stage1_c45_s_fa3), .Co(stage1_c45_c_fa3));
    FA fa_329(.A(stage0_r17_c28), .B(stage0_r18_c27), .C(stage0_r19_c26), .So(stage1_c45_s_fa4), .Co(stage1_c45_c_fa4));
    FA fa_330(.A(stage0_r20_c25), .B(stage0_r21_c24), .C(stage0_r22_c23), .So(stage1_c45_s_fa5), .Co(stage1_c45_c_fa5));
    FA fa_331(.A(stage0_r23_c22), .B(stage0_r24_c21), .C(stage0_r25_c20), .So(stage1_c45_s_fa6), .Co(stage1_c45_c_fa6));
    FA fa_332(.A(stage0_r26_c19), .B(stage0_r27_c18), .C(stage0_r28_c17), .So(stage1_c45_s_fa7), .Co(stage1_c45_c_fa7));
    FA fa_333(.A(stage0_r29_c16), .B(stage0_r30_c15), .C(stage0_r31_c14), .So(stage1_c45_s_fa8), .Co(stage1_c45_c_fa8));
    FA fa_334(.A(stage0_r32_c13), .B(stage0_r33_c12), .C(stage0_r34_c11), .So(stage1_c45_s_fa9), .Co(stage1_c45_c_fa9));
    FA fa_335(.A(stage0_r35_c10), .B(stage0_r36_c9), .C(stage0_r37_c8), .So(stage1_c45_s_fa10), .Co(stage1_c45_c_fa10));
    FA fa_336(.A(stage0_r38_c7), .B(stage0_r39_c6), .C(stage0_r40_c5), .So(stage1_c45_s_fa11), .Co(stage1_c45_c_fa11));
    FA fa_337(.A(stage0_r41_c4), .B(stage0_r42_c3), .C(stage0_r43_c2), .So(stage1_c45_s_fa12), .Co(stage1_c45_c_fa12));
    HA ha_18(.A(stage0_r44_c1), .B(stage0_r45_c0), .So(stage1_c45_s_ha0), .Co(stage1_c45_c_ha0));
    FA fa_338(.A(stage0_r6_c40), .B(stage0_r7_c39), .C(stage0_r8_c38), .So(stage1_c46_s_fa0), .Co(stage1_c46_c_fa0));
    FA fa_339(.A(stage0_r9_c37), .B(stage0_r10_c36), .C(stage0_r11_c35), .So(stage1_c46_s_fa1), .Co(stage1_c46_c_fa1));
    FA fa_340(.A(stage0_r12_c34), .B(stage0_r13_c33), .C(stage0_r14_c32), .So(stage1_c46_s_fa2), .Co(stage1_c46_c_fa2));
    FA fa_341(.A(stage0_r15_c31), .B(stage0_r16_c30), .C(stage0_r17_c29), .So(stage1_c46_s_fa3), .Co(stage1_c46_c_fa3));
    FA fa_342(.A(stage0_r18_c28), .B(stage0_r19_c27), .C(stage0_r20_c26), .So(stage1_c46_s_fa4), .Co(stage1_c46_c_fa4));
    FA fa_343(.A(stage0_r21_c25), .B(stage0_r22_c24), .C(stage0_r23_c23), .So(stage1_c46_s_fa5), .Co(stage1_c46_c_fa5));
    FA fa_344(.A(stage0_r24_c22), .B(stage0_r25_c21), .C(stage0_r26_c20), .So(stage1_c46_s_fa6), .Co(stage1_c46_c_fa6));
    FA fa_345(.A(stage0_r27_c19), .B(stage0_r28_c18), .C(stage0_r29_c17), .So(stage1_c46_s_fa7), .Co(stage1_c46_c_fa7));
    FA fa_346(.A(stage0_r30_c16), .B(stage0_r31_c15), .C(stage0_r32_c14), .So(stage1_c46_s_fa8), .Co(stage1_c46_c_fa8));
    FA fa_347(.A(stage0_r33_c13), .B(stage0_r34_c12), .C(stage0_r35_c11), .So(stage1_c46_s_fa9), .Co(stage1_c46_c_fa9));
    FA fa_348(.A(stage0_r36_c10), .B(stage0_r37_c9), .C(stage0_r38_c8), .So(stage1_c46_s_fa10), .Co(stage1_c46_c_fa10));
    FA fa_349(.A(stage0_r39_c7), .B(stage0_r40_c6), .C(stage0_r41_c5), .So(stage1_c46_s_fa11), .Co(stage1_c46_c_fa11));
    FA fa_350(.A(stage0_r42_c4), .B(stage0_r43_c3), .C(stage0_r44_c2), .So(stage1_c46_s_fa12), .Co(stage1_c46_c_fa12));
    HA ha_19(.A(stage0_r45_c1), .B(stage0_r46_c0), .So(stage1_c46_s_ha0), .Co(stage1_c46_c_ha0));
    FA fa_351(.A(stage0_r7_c40), .B(stage0_r8_c39), .C(stage0_r9_c38), .So(stage1_c47_s_fa0), .Co(stage1_c47_c_fa0));
    FA fa_352(.A(stage0_r10_c37), .B(stage0_r11_c36), .C(stage0_r12_c35), .So(stage1_c47_s_fa1), .Co(stage1_c47_c_fa1));
    FA fa_353(.A(stage0_r13_c34), .B(stage0_r14_c33), .C(stage0_r15_c32), .So(stage1_c47_s_fa2), .Co(stage1_c47_c_fa2));
    FA fa_354(.A(stage0_r16_c31), .B(stage0_r17_c30), .C(stage0_r18_c29), .So(stage1_c47_s_fa3), .Co(stage1_c47_c_fa3));
    FA fa_355(.A(stage0_r19_c28), .B(stage0_r20_c27), .C(stage0_r21_c26), .So(stage1_c47_s_fa4), .Co(stage1_c47_c_fa4));
    FA fa_356(.A(stage0_r22_c25), .B(stage0_r23_c24), .C(stage0_r24_c23), .So(stage1_c47_s_fa5), .Co(stage1_c47_c_fa5));
    FA fa_357(.A(stage0_r25_c22), .B(stage0_r26_c21), .C(stage0_r27_c20), .So(stage1_c47_s_fa6), .Co(stage1_c47_c_fa6));
    FA fa_358(.A(stage0_r28_c19), .B(stage0_r29_c18), .C(stage0_r30_c17), .So(stage1_c47_s_fa7), .Co(stage1_c47_c_fa7));
    FA fa_359(.A(stage0_r31_c16), .B(stage0_r32_c15), .C(stage0_r33_c14), .So(stage1_c47_s_fa8), .Co(stage1_c47_c_fa8));
    FA fa_360(.A(stage0_r34_c13), .B(stage0_r35_c12), .C(stage0_r36_c11), .So(stage1_c47_s_fa9), .Co(stage1_c47_c_fa9));
    FA fa_361(.A(stage0_r37_c10), .B(stage0_r38_c9), .C(stage0_r39_c8), .So(stage1_c47_s_fa10), .Co(stage1_c47_c_fa10));
    FA fa_362(.A(stage0_r40_c7), .B(stage0_r41_c6), .C(stage0_r42_c5), .So(stage1_c47_s_fa11), .Co(stage1_c47_c_fa11));
    FA fa_363(.A(stage0_r43_c4), .B(stage0_r44_c3), .C(stage0_r45_c2), .So(stage1_c47_s_fa12), .Co(stage1_c47_c_fa12));
    HA ha_20(.A(stage0_r46_c1), .B(stage0_r47_c0), .So(stage1_c47_s_ha0), .Co(stage1_c47_c_ha0));
    FA fa_364(.A(stage0_r8_c40), .B(stage0_r9_c39), .C(stage0_r10_c38), .So(stage1_c48_s_fa0), .Co(stage1_c48_c_fa0));
    FA fa_365(.A(stage0_r11_c37), .B(stage0_r12_c36), .C(stage0_r13_c35), .So(stage1_c48_s_fa1), .Co(stage1_c48_c_fa1));
    FA fa_366(.A(stage0_r14_c34), .B(stage0_r15_c33), .C(stage0_r16_c32), .So(stage1_c48_s_fa2), .Co(stage1_c48_c_fa2));
    FA fa_367(.A(stage0_r17_c31), .B(stage0_r18_c30), .C(stage0_r19_c29), .So(stage1_c48_s_fa3), .Co(stage1_c48_c_fa3));
    FA fa_368(.A(stage0_r20_c28), .B(stage0_r21_c27), .C(stage0_r22_c26), .So(stage1_c48_s_fa4), .Co(stage1_c48_c_fa4));
    FA fa_369(.A(stage0_r23_c25), .B(stage0_r24_c24), .C(stage0_r25_c23), .So(stage1_c48_s_fa5), .Co(stage1_c48_c_fa5));
    FA fa_370(.A(stage0_r26_c22), .B(stage0_r27_c21), .C(stage0_r28_c20), .So(stage1_c48_s_fa6), .Co(stage1_c48_c_fa6));
    FA fa_371(.A(stage0_r29_c19), .B(stage0_r30_c18), .C(stage0_r31_c17), .So(stage1_c48_s_fa7), .Co(stage1_c48_c_fa7));
    FA fa_372(.A(stage0_r32_c16), .B(stage0_r33_c15), .C(stage0_r34_c14), .So(stage1_c48_s_fa8), .Co(stage1_c48_c_fa8));
    FA fa_373(.A(stage0_r35_c13), .B(stage0_r36_c12), .C(stage0_r37_c11), .So(stage1_c48_s_fa9), .Co(stage1_c48_c_fa9));
    FA fa_374(.A(stage0_r38_c10), .B(stage0_r39_c9), .C(stage0_r40_c8), .So(stage1_c48_s_fa10), .Co(stage1_c48_c_fa10));
    FA fa_375(.A(stage0_r41_c7), .B(stage0_r42_c6), .C(stage0_r43_c5), .So(stage1_c48_s_fa11), .Co(stage1_c48_c_fa11));
    FA fa_376(.A(stage0_r44_c4), .B(stage0_r45_c3), .C(stage0_r46_c2), .So(stage1_c48_s_fa12), .Co(stage1_c48_c_fa12));
    HA ha_21(.A(stage0_r47_c1), .B(stage0_r48_c0), .So(stage1_c48_s_ha0), .Co(stage1_c48_c_ha0));
    FA fa_377(.A(stage0_r9_c40), .B(stage0_r10_c39), .C(stage0_r11_c38), .So(stage1_c49_s_fa0), .Co(stage1_c49_c_fa0));
    FA fa_378(.A(stage0_r12_c37), .B(stage0_r13_c36), .C(stage0_r14_c35), .So(stage1_c49_s_fa1), .Co(stage1_c49_c_fa1));
    FA fa_379(.A(stage0_r15_c34), .B(stage0_r16_c33), .C(stage0_r17_c32), .So(stage1_c49_s_fa2), .Co(stage1_c49_c_fa2));
    FA fa_380(.A(stage0_r18_c31), .B(stage0_r19_c30), .C(stage0_r20_c29), .So(stage1_c49_s_fa3), .Co(stage1_c49_c_fa3));
    FA fa_381(.A(stage0_r21_c28), .B(stage0_r22_c27), .C(stage0_r23_c26), .So(stage1_c49_s_fa4), .Co(stage1_c49_c_fa4));
    FA fa_382(.A(stage0_r24_c25), .B(stage0_r25_c24), .C(stage0_r26_c23), .So(stage1_c49_s_fa5), .Co(stage1_c49_c_fa5));
    FA fa_383(.A(stage0_r27_c22), .B(stage0_r28_c21), .C(stage0_r29_c20), .So(stage1_c49_s_fa6), .Co(stage1_c49_c_fa6));
    FA fa_384(.A(stage0_r30_c19), .B(stage0_r31_c18), .C(stage0_r32_c17), .So(stage1_c49_s_fa7), .Co(stage1_c49_c_fa7));
    FA fa_385(.A(stage0_r33_c16), .B(stage0_r34_c15), .C(stage0_r35_c14), .So(stage1_c49_s_fa8), .Co(stage1_c49_c_fa8));
    FA fa_386(.A(stage0_r36_c13), .B(stage0_r37_c12), .C(stage0_r38_c11), .So(stage1_c49_s_fa9), .Co(stage1_c49_c_fa9));
    FA fa_387(.A(stage0_r39_c10), .B(stage0_r40_c9), .C(stage0_r41_c8), .So(stage1_c49_s_fa10), .Co(stage1_c49_c_fa10));
    FA fa_388(.A(stage0_r42_c7), .B(stage0_r43_c6), .C(stage0_r44_c5), .So(stage1_c49_s_fa11), .Co(stage1_c49_c_fa11));
    FA fa_389(.A(stage0_r45_c4), .B(stage0_r46_c3), .C(stage0_r47_c2), .So(stage1_c49_s_fa12), .Co(stage1_c49_c_fa12));
    HA ha_22(.A(stage0_r48_c1), .B(stage0_r49_c0), .So(stage1_c49_s_ha0), .Co(stage1_c49_c_ha0));
    FA fa_390(.A(stage0_r10_c40), .B(stage0_r11_c39), .C(stage0_r12_c38), .So(stage1_c50_s_fa0), .Co(stage1_c50_c_fa0));
    FA fa_391(.A(stage0_r13_c37), .B(stage0_r14_c36), .C(stage0_r15_c35), .So(stage1_c50_s_fa1), .Co(stage1_c50_c_fa1));
    FA fa_392(.A(stage0_r16_c34), .B(stage0_r17_c33), .C(stage0_r18_c32), .So(stage1_c50_s_fa2), .Co(stage1_c50_c_fa2));
    FA fa_393(.A(stage0_r19_c31), .B(stage0_r20_c30), .C(stage0_r21_c29), .So(stage1_c50_s_fa3), .Co(stage1_c50_c_fa3));
    FA fa_394(.A(stage0_r22_c28), .B(stage0_r23_c27), .C(stage0_r24_c26), .So(stage1_c50_s_fa4), .Co(stage1_c50_c_fa4));
    FA fa_395(.A(stage0_r25_c25), .B(stage0_r26_c24), .C(stage0_r27_c23), .So(stage1_c50_s_fa5), .Co(stage1_c50_c_fa5));
    FA fa_396(.A(stage0_r28_c22), .B(stage0_r29_c21), .C(stage0_r30_c20), .So(stage1_c50_s_fa6), .Co(stage1_c50_c_fa6));
    FA fa_397(.A(stage0_r31_c19), .B(stage0_r32_c18), .C(stage0_r33_c17), .So(stage1_c50_s_fa7), .Co(stage1_c50_c_fa7));
    FA fa_398(.A(stage0_r34_c16), .B(stage0_r35_c15), .C(stage0_r36_c14), .So(stage1_c50_s_fa8), .Co(stage1_c50_c_fa8));
    FA fa_399(.A(stage0_r37_c13), .B(stage0_r38_c12), .C(stage0_r39_c11), .So(stage1_c50_s_fa9), .Co(stage1_c50_c_fa9));
    FA fa_400(.A(stage0_r40_c10), .B(stage0_r41_c9), .C(stage0_r42_c8), .So(stage1_c50_s_fa10), .Co(stage1_c50_c_fa10));
    FA fa_401(.A(stage0_r43_c7), .B(stage0_r44_c6), .C(stage0_r45_c5), .So(stage1_c50_s_fa11), .Co(stage1_c50_c_fa11));
    FA fa_402(.A(stage0_r46_c4), .B(stage0_r47_c3), .C(stage0_r48_c2), .So(stage1_c50_s_fa12), .Co(stage1_c50_c_fa12));
    HA ha_23(.A(stage0_r49_c1), .B(stage0_r50_c0), .So(stage1_c50_s_ha0), .Co(stage1_c50_c_ha0));
    FA fa_403(.A(stage0_r11_c40), .B(stage0_r12_c39), .C(stage0_r13_c38), .So(stage1_c51_s_fa0), .Co(stage1_c51_c_fa0));
    FA fa_404(.A(stage0_r14_c37), .B(stage0_r15_c36), .C(stage0_r16_c35), .So(stage1_c51_s_fa1), .Co(stage1_c51_c_fa1));
    FA fa_405(.A(stage0_r17_c34), .B(stage0_r18_c33), .C(stage0_r19_c32), .So(stage1_c51_s_fa2), .Co(stage1_c51_c_fa2));
    FA fa_406(.A(stage0_r20_c31), .B(stage0_r21_c30), .C(stage0_r22_c29), .So(stage1_c51_s_fa3), .Co(stage1_c51_c_fa3));
    FA fa_407(.A(stage0_r23_c28), .B(stage0_r24_c27), .C(stage0_r25_c26), .So(stage1_c51_s_fa4), .Co(stage1_c51_c_fa4));
    FA fa_408(.A(stage0_r26_c25), .B(stage0_r27_c24), .C(stage0_r28_c23), .So(stage1_c51_s_fa5), .Co(stage1_c51_c_fa5));
    FA fa_409(.A(stage0_r29_c22), .B(stage0_r30_c21), .C(stage0_r31_c20), .So(stage1_c51_s_fa6), .Co(stage1_c51_c_fa6));
    FA fa_410(.A(stage0_r32_c19), .B(stage0_r33_c18), .C(stage0_r34_c17), .So(stage1_c51_s_fa7), .Co(stage1_c51_c_fa7));
    FA fa_411(.A(stage0_r35_c16), .B(stage0_r36_c15), .C(stage0_r37_c14), .So(stage1_c51_s_fa8), .Co(stage1_c51_c_fa8));
    FA fa_412(.A(stage0_r38_c13), .B(stage0_r39_c12), .C(stage0_r40_c11), .So(stage1_c51_s_fa9), .Co(stage1_c51_c_fa9));
    FA fa_413(.A(stage0_r41_c10), .B(stage0_r42_c9), .C(stage0_r43_c8), .So(stage1_c51_s_fa10), .Co(stage1_c51_c_fa10));
    FA fa_414(.A(stage0_r44_c7), .B(stage0_r45_c6), .C(stage0_r46_c5), .So(stage1_c51_s_fa11), .Co(stage1_c51_c_fa11));
    FA fa_415(.A(stage0_r47_c4), .B(stage0_r48_c3), .C(stage0_r49_c2), .So(stage1_c51_s_fa12), .Co(stage1_c51_c_fa12));
    HA ha_24(.A(stage0_r50_c1), .B(stage0_r51_c0), .So(stage1_c51_s_ha0), .Co(stage1_c51_c_ha0));
    FA fa_416(.A(stage0_r12_c40), .B(stage0_r13_c39), .C(stage0_r14_c38), .So(stage1_c52_s_fa0), .Co(stage1_c52_c_fa0));
    FA fa_417(.A(stage0_r15_c37), .B(stage0_r16_c36), .C(stage0_r17_c35), .So(stage1_c52_s_fa1), .Co(stage1_c52_c_fa1));
    FA fa_418(.A(stage0_r18_c34), .B(stage0_r19_c33), .C(stage0_r20_c32), .So(stage1_c52_s_fa2), .Co(stage1_c52_c_fa2));
    FA fa_419(.A(stage0_r21_c31), .B(stage0_r22_c30), .C(stage0_r23_c29), .So(stage1_c52_s_fa3), .Co(stage1_c52_c_fa3));
    FA fa_420(.A(stage0_r24_c28), .B(stage0_r25_c27), .C(stage0_r26_c26), .So(stage1_c52_s_fa4), .Co(stage1_c52_c_fa4));
    FA fa_421(.A(stage0_r27_c25), .B(stage0_r28_c24), .C(stage0_r29_c23), .So(stage1_c52_s_fa5), .Co(stage1_c52_c_fa5));
    FA fa_422(.A(stage0_r30_c22), .B(stage0_r31_c21), .C(stage0_r32_c20), .So(stage1_c52_s_fa6), .Co(stage1_c52_c_fa6));
    FA fa_423(.A(stage0_r33_c19), .B(stage0_r34_c18), .C(stage0_r35_c17), .So(stage1_c52_s_fa7), .Co(stage1_c52_c_fa7));
    FA fa_424(.A(stage0_r36_c16), .B(stage0_r37_c15), .C(stage0_r38_c14), .So(stage1_c52_s_fa8), .Co(stage1_c52_c_fa8));
    FA fa_425(.A(stage0_r39_c13), .B(stage0_r40_c12), .C(stage0_r41_c11), .So(stage1_c52_s_fa9), .Co(stage1_c52_c_fa9));
    FA fa_426(.A(stage0_r42_c10), .B(stage0_r43_c9), .C(stage0_r44_c8), .So(stage1_c52_s_fa10), .Co(stage1_c52_c_fa10));
    FA fa_427(.A(stage0_r45_c7), .B(stage0_r46_c6), .C(stage0_r47_c5), .So(stage1_c52_s_fa11), .Co(stage1_c52_c_fa11));
    FA fa_428(.A(stage0_r48_c4), .B(stage0_r49_c3), .C(stage0_r50_c2), .So(stage1_c52_s_fa12), .Co(stage1_c52_c_fa12));
    HA ha_25(.A(stage0_r51_c1), .B(stage0_r52_c0), .So(stage1_c52_s_ha0), .Co(stage1_c52_c_ha0));
    FA fa_429(.A(stage0_r13_c40), .B(stage0_r14_c39), .C(stage0_r15_c38), .So(stage1_c53_s_fa0), .Co(stage1_c53_c_fa0));
    FA fa_430(.A(stage0_r16_c37), .B(stage0_r17_c36), .C(stage0_r18_c35), .So(stage1_c53_s_fa1), .Co(stage1_c53_c_fa1));
    FA fa_431(.A(stage0_r19_c34), .B(stage0_r20_c33), .C(stage0_r21_c32), .So(stage1_c53_s_fa2), .Co(stage1_c53_c_fa2));
    FA fa_432(.A(stage0_r22_c31), .B(stage0_r23_c30), .C(stage0_r24_c29), .So(stage1_c53_s_fa3), .Co(stage1_c53_c_fa3));
    FA fa_433(.A(stage0_r25_c28), .B(stage0_r26_c27), .C(stage0_r27_c26), .So(stage1_c53_s_fa4), .Co(stage1_c53_c_fa4));
    FA fa_434(.A(stage0_r28_c25), .B(stage0_r29_c24), .C(stage0_r30_c23), .So(stage1_c53_s_fa5), .Co(stage1_c53_c_fa5));
    FA fa_435(.A(stage0_r31_c22), .B(stage0_r32_c21), .C(stage0_r33_c20), .So(stage1_c53_s_fa6), .Co(stage1_c53_c_fa6));
    FA fa_436(.A(stage0_r34_c19), .B(stage0_r35_c18), .C(stage0_r36_c17), .So(stage1_c53_s_fa7), .Co(stage1_c53_c_fa7));
    FA fa_437(.A(stage0_r37_c16), .B(stage0_r38_c15), .C(stage0_r39_c14), .So(stage1_c53_s_fa8), .Co(stage1_c53_c_fa8));
    FA fa_438(.A(stage0_r40_c13), .B(stage0_r41_c12), .C(stage0_r42_c11), .So(stage1_c53_s_fa9), .Co(stage1_c53_c_fa9));
    FA fa_439(.A(stage0_r43_c10), .B(stage0_r44_c9), .C(stage0_r45_c8), .So(stage1_c53_s_fa10), .Co(stage1_c53_c_fa10));
    FA fa_440(.A(stage0_r46_c7), .B(stage0_r47_c6), .C(stage0_r48_c5), .So(stage1_c53_s_fa11), .Co(stage1_c53_c_fa11));
    FA fa_441(.A(stage0_r49_c4), .B(stage0_r50_c3), .C(stage0_r51_c2), .So(stage1_c53_s_fa12), .Co(stage1_c53_c_fa12));
    HA ha_26(.A(stage0_r52_c1), .B(stage0_r53_c0), .So(stage1_c53_s_ha0), .Co(stage1_c53_c_ha0));
    FA fa_442(.A(stage0_r14_c40), .B(stage0_r15_c39), .C(stage0_r16_c38), .So(stage1_c54_s_fa0), .Co(stage1_c54_c_fa0));
    FA fa_443(.A(stage0_r17_c37), .B(stage0_r18_c36), .C(stage0_r19_c35), .So(stage1_c54_s_fa1), .Co(stage1_c54_c_fa1));
    FA fa_444(.A(stage0_r20_c34), .B(stage0_r21_c33), .C(stage0_r22_c32), .So(stage1_c54_s_fa2), .Co(stage1_c54_c_fa2));
    FA fa_445(.A(stage0_r23_c31), .B(stage0_r24_c30), .C(stage0_r25_c29), .So(stage1_c54_s_fa3), .Co(stage1_c54_c_fa3));
    FA fa_446(.A(stage0_r26_c28), .B(stage0_r27_c27), .C(stage0_r28_c26), .So(stage1_c54_s_fa4), .Co(stage1_c54_c_fa4));
    FA fa_447(.A(stage0_r29_c25), .B(stage0_r30_c24), .C(stage0_r31_c23), .So(stage1_c54_s_fa5), .Co(stage1_c54_c_fa5));
    FA fa_448(.A(stage0_r32_c22), .B(stage0_r33_c21), .C(stage0_r34_c20), .So(stage1_c54_s_fa6), .Co(stage1_c54_c_fa6));
    FA fa_449(.A(stage0_r35_c19), .B(stage0_r36_c18), .C(stage0_r37_c17), .So(stage1_c54_s_fa7), .Co(stage1_c54_c_fa7));
    FA fa_450(.A(stage0_r38_c16), .B(stage0_r39_c15), .C(stage0_r40_c14), .So(stage1_c54_s_fa8), .Co(stage1_c54_c_fa8));
    FA fa_451(.A(stage0_r41_c13), .B(stage0_r42_c12), .C(stage0_r43_c11), .So(stage1_c54_s_fa9), .Co(stage1_c54_c_fa9));
    FA fa_452(.A(stage0_r44_c10), .B(stage0_r45_c9), .C(stage0_r46_c8), .So(stage1_c54_s_fa10), .Co(stage1_c54_c_fa10));
    FA fa_453(.A(stage0_r47_c7), .B(stage0_r48_c6), .C(stage0_r49_c5), .So(stage1_c54_s_fa11), .Co(stage1_c54_c_fa11));
    FA fa_454(.A(stage0_r50_c4), .B(stage0_r51_c3), .C(stage0_r52_c2), .So(stage1_c54_s_fa12), .Co(stage1_c54_c_fa12));
    HA ha_27(.A(stage0_r53_c1), .B(stage0_r54_c0), .So(stage1_c54_s_ha0), .Co(stage1_c54_c_ha0));
    FA fa_455(.A(stage0_r15_c40), .B(stage0_r16_c39), .C(stage0_r17_c38), .So(stage1_c55_s_fa0), .Co(stage1_c55_c_fa0));
    FA fa_456(.A(stage0_r18_c37), .B(stage0_r19_c36), .C(stage0_r20_c35), .So(stage1_c55_s_fa1), .Co(stage1_c55_c_fa1));
    FA fa_457(.A(stage0_r21_c34), .B(stage0_r22_c33), .C(stage0_r23_c32), .So(stage1_c55_s_fa2), .Co(stage1_c55_c_fa2));
    FA fa_458(.A(stage0_r24_c31), .B(stage0_r25_c30), .C(stage0_r26_c29), .So(stage1_c55_s_fa3), .Co(stage1_c55_c_fa3));
    FA fa_459(.A(stage0_r27_c28), .B(stage0_r28_c27), .C(stage0_r29_c26), .So(stage1_c55_s_fa4), .Co(stage1_c55_c_fa4));
    FA fa_460(.A(stage0_r30_c25), .B(stage0_r31_c24), .C(stage0_r32_c23), .So(stage1_c55_s_fa5), .Co(stage1_c55_c_fa5));
    FA fa_461(.A(stage0_r33_c22), .B(stage0_r34_c21), .C(stage0_r35_c20), .So(stage1_c55_s_fa6), .Co(stage1_c55_c_fa6));
    FA fa_462(.A(stage0_r36_c19), .B(stage0_r37_c18), .C(stage0_r38_c17), .So(stage1_c55_s_fa7), .Co(stage1_c55_c_fa7));
    FA fa_463(.A(stage0_r39_c16), .B(stage0_r40_c15), .C(stage0_r41_c14), .So(stage1_c55_s_fa8), .Co(stage1_c55_c_fa8));
    FA fa_464(.A(stage0_r42_c13), .B(stage0_r43_c12), .C(stage0_r44_c11), .So(stage1_c55_s_fa9), .Co(stage1_c55_c_fa9));
    FA fa_465(.A(stage0_r45_c10), .B(stage0_r46_c9), .C(stage0_r47_c8), .So(stage1_c55_s_fa10), .Co(stage1_c55_c_fa10));
    FA fa_466(.A(stage0_r48_c7), .B(stage0_r49_c6), .C(stage0_r50_c5), .So(stage1_c55_s_fa11), .Co(stage1_c55_c_fa11));
    FA fa_467(.A(stage0_r51_c4), .B(stage0_r52_c3), .C(stage0_r53_c2), .So(stage1_c55_s_fa12), .Co(stage1_c55_c_fa12));
    HA ha_28(.A(stage0_r54_c1), .B(stage0_r55_c0), .So(stage1_c55_s_ha0), .Co(stage1_c55_c_ha0));
    FA fa_468(.A(stage0_r16_c40), .B(stage0_r17_c39), .C(stage0_r18_c38), .So(stage1_c56_s_fa0), .Co(stage1_c56_c_fa0));
    FA fa_469(.A(stage0_r19_c37), .B(stage0_r20_c36), .C(stage0_r21_c35), .So(stage1_c56_s_fa1), .Co(stage1_c56_c_fa1));
    FA fa_470(.A(stage0_r22_c34), .B(stage0_r23_c33), .C(stage0_r24_c32), .So(stage1_c56_s_fa2), .Co(stage1_c56_c_fa2));
    FA fa_471(.A(stage0_r25_c31), .B(stage0_r26_c30), .C(stage0_r27_c29), .So(stage1_c56_s_fa3), .Co(stage1_c56_c_fa3));
    FA fa_472(.A(stage0_r28_c28), .B(stage0_r29_c27), .C(stage0_r30_c26), .So(stage1_c56_s_fa4), .Co(stage1_c56_c_fa4));
    FA fa_473(.A(stage0_r31_c25), .B(stage0_r32_c24), .C(stage0_r33_c23), .So(stage1_c56_s_fa5), .Co(stage1_c56_c_fa5));
    FA fa_474(.A(stage0_r34_c22), .B(stage0_r35_c21), .C(stage0_r36_c20), .So(stage1_c56_s_fa6), .Co(stage1_c56_c_fa6));
    FA fa_475(.A(stage0_r37_c19), .B(stage0_r38_c18), .C(stage0_r39_c17), .So(stage1_c56_s_fa7), .Co(stage1_c56_c_fa7));
    FA fa_476(.A(stage0_r40_c16), .B(stage0_r41_c15), .C(stage0_r42_c14), .So(stage1_c56_s_fa8), .Co(stage1_c56_c_fa8));
    FA fa_477(.A(stage0_r43_c13), .B(stage0_r44_c12), .C(stage0_r45_c11), .So(stage1_c56_s_fa9), .Co(stage1_c56_c_fa9));
    FA fa_478(.A(stage0_r46_c10), .B(stage0_r47_c9), .C(stage0_r48_c8), .So(stage1_c56_s_fa10), .Co(stage1_c56_c_fa10));
    FA fa_479(.A(stage0_r49_c7), .B(stage0_r50_c6), .C(stage0_r51_c5), .So(stage1_c56_s_fa11), .Co(stage1_c56_c_fa11));
    FA fa_480(.A(stage0_r52_c4), .B(stage0_r53_c3), .C(stage0_r54_c2), .So(stage1_c56_s_fa12), .Co(stage1_c56_c_fa12));
    HA ha_29(.A(stage0_r55_c1), .B(stage0_r56_c0), .So(stage1_c56_s_ha0), .Co(stage1_c56_c_ha0));
    FA fa_481(.A(stage0_r17_c40), .B(stage0_r18_c39), .C(stage0_r19_c38), .So(stage1_c57_s_fa0), .Co(stage1_c57_c_fa0));
    FA fa_482(.A(stage0_r20_c37), .B(stage0_r21_c36), .C(stage0_r22_c35), .So(stage1_c57_s_fa1), .Co(stage1_c57_c_fa1));
    FA fa_483(.A(stage0_r23_c34), .B(stage0_r24_c33), .C(stage0_r25_c32), .So(stage1_c57_s_fa2), .Co(stage1_c57_c_fa2));
    FA fa_484(.A(stage0_r26_c31), .B(stage0_r27_c30), .C(stage0_r28_c29), .So(stage1_c57_s_fa3), .Co(stage1_c57_c_fa3));
    FA fa_485(.A(stage0_r29_c28), .B(stage0_r30_c27), .C(stage0_r31_c26), .So(stage1_c57_s_fa4), .Co(stage1_c57_c_fa4));
    FA fa_486(.A(stage0_r32_c25), .B(stage0_r33_c24), .C(stage0_r34_c23), .So(stage1_c57_s_fa5), .Co(stage1_c57_c_fa5));
    FA fa_487(.A(stage0_r35_c22), .B(stage0_r36_c21), .C(stage0_r37_c20), .So(stage1_c57_s_fa6), .Co(stage1_c57_c_fa6));
    FA fa_488(.A(stage0_r38_c19), .B(stage0_r39_c18), .C(stage0_r40_c17), .So(stage1_c57_s_fa7), .Co(stage1_c57_c_fa7));
    FA fa_489(.A(stage0_r41_c16), .B(stage0_r42_c15), .C(stage0_r43_c14), .So(stage1_c57_s_fa8), .Co(stage1_c57_c_fa8));
    FA fa_490(.A(stage0_r44_c13), .B(stage0_r45_c12), .C(stage0_r46_c11), .So(stage1_c57_s_fa9), .Co(stage1_c57_c_fa9));
    FA fa_491(.A(stage0_r47_c10), .B(stage0_r48_c9), .C(stage0_r49_c8), .So(stage1_c57_s_fa10), .Co(stage1_c57_c_fa10));
    FA fa_492(.A(stage0_r50_c7), .B(stage0_r51_c6), .C(stage0_r52_c5), .So(stage1_c57_s_fa11), .Co(stage1_c57_c_fa11));
    FA fa_493(.A(stage0_r53_c4), .B(stage0_r54_c3), .C(stage0_r55_c2), .So(stage1_c57_s_fa12), .Co(stage1_c57_c_fa12));
    HA ha_30(.A(stage0_r56_c1), .B(stage0_r57_c0), .So(stage1_c57_s_ha0), .Co(stage1_c57_c_ha0));
    FA fa_494(.A(stage0_r18_c40), .B(stage0_r19_c39), .C(stage0_r20_c38), .So(stage1_c58_s_fa0), .Co(stage1_c58_c_fa0));
    FA fa_495(.A(stage0_r21_c37), .B(stage0_r22_c36), .C(stage0_r23_c35), .So(stage1_c58_s_fa1), .Co(stage1_c58_c_fa1));
    FA fa_496(.A(stage0_r24_c34), .B(stage0_r25_c33), .C(stage0_r26_c32), .So(stage1_c58_s_fa2), .Co(stage1_c58_c_fa2));
    FA fa_497(.A(stage0_r27_c31), .B(stage0_r28_c30), .C(stage0_r29_c29), .So(stage1_c58_s_fa3), .Co(stage1_c58_c_fa3));
    FA fa_498(.A(stage0_r30_c28), .B(stage0_r31_c27), .C(stage0_r32_c26), .So(stage1_c58_s_fa4), .Co(stage1_c58_c_fa4));
    FA fa_499(.A(stage0_r33_c25), .B(stage0_r34_c24), .C(stage0_r35_c23), .So(stage1_c58_s_fa5), .Co(stage1_c58_c_fa5));
    FA fa_500(.A(stage0_r36_c22), .B(stage0_r37_c21), .C(stage0_r38_c20), .So(stage1_c58_s_fa6), .Co(stage1_c58_c_fa6));
    FA fa_501(.A(stage0_r39_c19), .B(stage0_r40_c18), .C(stage0_r41_c17), .So(stage1_c58_s_fa7), .Co(stage1_c58_c_fa7));
    FA fa_502(.A(stage0_r42_c16), .B(stage0_r43_c15), .C(stage0_r44_c14), .So(stage1_c58_s_fa8), .Co(stage1_c58_c_fa8));
    FA fa_503(.A(stage0_r45_c13), .B(stage0_r46_c12), .C(stage0_r47_c11), .So(stage1_c58_s_fa9), .Co(stage1_c58_c_fa9));
    FA fa_504(.A(stage0_r48_c10), .B(stage0_r49_c9), .C(stage0_r50_c8), .So(stage1_c58_s_fa10), .Co(stage1_c58_c_fa10));
    FA fa_505(.A(stage0_r51_c7), .B(stage0_r52_c6), .C(stage0_r53_c5), .So(stage1_c58_s_fa11), .Co(stage1_c58_c_fa11));
    FA fa_506(.A(stage0_r54_c4), .B(stage0_r55_c3), .C(stage0_r56_c2), .So(stage1_c58_s_fa12), .Co(stage1_c58_c_fa12));
    HA ha_31(.A(stage0_r57_c1), .B(stage0_r58_c0), .So(stage1_c58_s_ha0), .Co(stage1_c58_c_ha0));
    FA fa_507(.A(stage0_r19_c40), .B(stage0_r20_c39), .C(stage0_r21_c38), .So(stage1_c59_s_fa0), .Co(stage1_c59_c_fa0));
    FA fa_508(.A(stage0_r22_c37), .B(stage0_r23_c36), .C(stage0_r24_c35), .So(stage1_c59_s_fa1), .Co(stage1_c59_c_fa1));
    FA fa_509(.A(stage0_r25_c34), .B(stage0_r26_c33), .C(stage0_r27_c32), .So(stage1_c59_s_fa2), .Co(stage1_c59_c_fa2));
    FA fa_510(.A(stage0_r28_c31), .B(stage0_r29_c30), .C(stage0_r30_c29), .So(stage1_c59_s_fa3), .Co(stage1_c59_c_fa3));
    FA fa_511(.A(stage0_r31_c28), .B(stage0_r32_c27), .C(stage0_r33_c26), .So(stage1_c59_s_fa4), .Co(stage1_c59_c_fa4));
    FA fa_512(.A(stage0_r34_c25), .B(stage0_r35_c24), .C(stage0_r36_c23), .So(stage1_c59_s_fa5), .Co(stage1_c59_c_fa5));
    FA fa_513(.A(stage0_r37_c22), .B(stage0_r38_c21), .C(stage0_r39_c20), .So(stage1_c59_s_fa6), .Co(stage1_c59_c_fa6));
    FA fa_514(.A(stage0_r40_c19), .B(stage0_r41_c18), .C(stage0_r42_c17), .So(stage1_c59_s_fa7), .Co(stage1_c59_c_fa7));
    FA fa_515(.A(stage0_r43_c16), .B(stage0_r44_c15), .C(stage0_r45_c14), .So(stage1_c59_s_fa8), .Co(stage1_c59_c_fa8));
    FA fa_516(.A(stage0_r46_c13), .B(stage0_r47_c12), .C(stage0_r48_c11), .So(stage1_c59_s_fa9), .Co(stage1_c59_c_fa9));
    FA fa_517(.A(stage0_r49_c10), .B(stage0_r50_c9), .C(stage0_r51_c8), .So(stage1_c59_s_fa10), .Co(stage1_c59_c_fa10));
    FA fa_518(.A(stage0_r52_c7), .B(stage0_r53_c6), .C(stage0_r54_c5), .So(stage1_c59_s_fa11), .Co(stage1_c59_c_fa11));
    FA fa_519(.A(stage0_r55_c4), .B(stage0_r56_c3), .C(stage0_r57_c2), .So(stage1_c59_s_fa12), .Co(stage1_c59_c_fa12));
    HA ha_32(.A(stage0_r58_c1), .B(stage0_r59_c0), .So(stage1_c59_s_ha0), .Co(stage1_c59_c_ha0));
    FA fa_520(.A(stage0_r20_c40), .B(stage0_r21_c39), .C(stage0_r22_c38), .So(stage1_c60_s_fa0), .Co(stage1_c60_c_fa0));
    FA fa_521(.A(stage0_r23_c37), .B(stage0_r24_c36), .C(stage0_r25_c35), .So(stage1_c60_s_fa1), .Co(stage1_c60_c_fa1));
    FA fa_522(.A(stage0_r26_c34), .B(stage0_r27_c33), .C(stage0_r28_c32), .So(stage1_c60_s_fa2), .Co(stage1_c60_c_fa2));
    FA fa_523(.A(stage0_r29_c31), .B(stage0_r30_c30), .C(stage0_r31_c29), .So(stage1_c60_s_fa3), .Co(stage1_c60_c_fa3));
    FA fa_524(.A(stage0_r32_c28), .B(stage0_r33_c27), .C(stage0_r34_c26), .So(stage1_c60_s_fa4), .Co(stage1_c60_c_fa4));
    FA fa_525(.A(stage0_r35_c25), .B(stage0_r36_c24), .C(stage0_r37_c23), .So(stage1_c60_s_fa5), .Co(stage1_c60_c_fa5));
    FA fa_526(.A(stage0_r38_c22), .B(stage0_r39_c21), .C(stage0_r40_c20), .So(stage1_c60_s_fa6), .Co(stage1_c60_c_fa6));
    FA fa_527(.A(stage0_r41_c19), .B(stage0_r42_c18), .C(stage0_r43_c17), .So(stage1_c60_s_fa7), .Co(stage1_c60_c_fa7));
    FA fa_528(.A(stage0_r44_c16), .B(stage0_r45_c15), .C(stage0_r46_c14), .So(stage1_c60_s_fa8), .Co(stage1_c60_c_fa8));
    FA fa_529(.A(stage0_r47_c13), .B(stage0_r48_c12), .C(stage0_r49_c11), .So(stage1_c60_s_fa9), .Co(stage1_c60_c_fa9));
    FA fa_530(.A(stage0_r50_c10), .B(stage0_r51_c9), .C(stage0_r52_c8), .So(stage1_c60_s_fa10), .Co(stage1_c60_c_fa10));
    FA fa_531(.A(stage0_r53_c7), .B(stage0_r54_c6), .C(stage0_r55_c5), .So(stage1_c60_s_fa11), .Co(stage1_c60_c_fa11));
    FA fa_532(.A(stage0_r56_c4), .B(stage0_r57_c3), .C(stage0_r58_c2), .So(stage1_c60_s_fa12), .Co(stage1_c60_c_fa12));
    HA ha_33(.A(stage0_r59_c1), .B(stage0_r60_c0), .So(stage1_c60_s_ha0), .Co(stage1_c60_c_ha0));
    FA fa_533(.A(stage0_r21_c40), .B(stage0_r22_c39), .C(stage0_r23_c38), .So(stage1_c61_s_fa0), .Co(stage1_c61_c_fa0));
    FA fa_534(.A(stage0_r24_c37), .B(stage0_r25_c36), .C(stage0_r26_c35), .So(stage1_c61_s_fa1), .Co(stage1_c61_c_fa1));
    FA fa_535(.A(stage0_r27_c34), .B(stage0_r28_c33), .C(stage0_r29_c32), .So(stage1_c61_s_fa2), .Co(stage1_c61_c_fa2));
    FA fa_536(.A(stage0_r30_c31), .B(stage0_r31_c30), .C(stage0_r32_c29), .So(stage1_c61_s_fa3), .Co(stage1_c61_c_fa3));
    FA fa_537(.A(stage0_r33_c28), .B(stage0_r34_c27), .C(stage0_r35_c26), .So(stage1_c61_s_fa4), .Co(stage1_c61_c_fa4));
    FA fa_538(.A(stage0_r36_c25), .B(stage0_r37_c24), .C(stage0_r38_c23), .So(stage1_c61_s_fa5), .Co(stage1_c61_c_fa5));
    FA fa_539(.A(stage0_r39_c22), .B(stage0_r40_c21), .C(stage0_r41_c20), .So(stage1_c61_s_fa6), .Co(stage1_c61_c_fa6));
    FA fa_540(.A(stage0_r42_c19), .B(stage0_r43_c18), .C(stage0_r44_c17), .So(stage1_c61_s_fa7), .Co(stage1_c61_c_fa7));
    FA fa_541(.A(stage0_r45_c16), .B(stage0_r46_c15), .C(stage0_r47_c14), .So(stage1_c61_s_fa8), .Co(stage1_c61_c_fa8));
    FA fa_542(.A(stage0_r48_c13), .B(stage0_r49_c12), .C(stage0_r50_c11), .So(stage1_c61_s_fa9), .Co(stage1_c61_c_fa9));
    FA fa_543(.A(stage0_r51_c10), .B(stage0_r52_c9), .C(stage0_r53_c8), .So(stage1_c61_s_fa10), .Co(stage1_c61_c_fa10));
    FA fa_544(.A(stage0_r54_c7), .B(stage0_r55_c6), .C(stage0_r56_c5), .So(stage1_c61_s_fa11), .Co(stage1_c61_c_fa11));
    FA fa_545(.A(stage0_r57_c4), .B(stage0_r58_c3), .C(stage0_r59_c2), .So(stage1_c61_s_fa12), .Co(stage1_c61_c_fa12));
    HA ha_34(.A(stage0_r60_c1), .B(stage0_r61_c0), .So(stage1_c61_s_ha0), .Co(stage1_c61_c_ha0));
    FA fa_546(.A(stage0_r22_c40), .B(stage0_r23_c39), .C(stage0_r24_c38), .So(stage1_c62_s_fa0), .Co(stage1_c62_c_fa0));
    FA fa_547(.A(stage0_r25_c37), .B(stage0_r26_c36), .C(stage0_r27_c35), .So(stage1_c62_s_fa1), .Co(stage1_c62_c_fa1));
    FA fa_548(.A(stage0_r28_c34), .B(stage0_r29_c33), .C(stage0_r30_c32), .So(stage1_c62_s_fa2), .Co(stage1_c62_c_fa2));
    FA fa_549(.A(stage0_r31_c31), .B(stage0_r32_c30), .C(stage0_r33_c29), .So(stage1_c62_s_fa3), .Co(stage1_c62_c_fa3));
    FA fa_550(.A(stage0_r34_c28), .B(stage0_r35_c27), .C(stage0_r36_c26), .So(stage1_c62_s_fa4), .Co(stage1_c62_c_fa4));
    FA fa_551(.A(stage0_r37_c25), .B(stage0_r38_c24), .C(stage0_r39_c23), .So(stage1_c62_s_fa5), .Co(stage1_c62_c_fa5));
    FA fa_552(.A(stage0_r40_c22), .B(stage0_r41_c21), .C(stage0_r42_c20), .So(stage1_c62_s_fa6), .Co(stage1_c62_c_fa6));
    FA fa_553(.A(stage0_r43_c19), .B(stage0_r44_c18), .C(stage0_r45_c17), .So(stage1_c62_s_fa7), .Co(stage1_c62_c_fa7));
    FA fa_554(.A(stage0_r46_c16), .B(stage0_r47_c15), .C(stage0_r48_c14), .So(stage1_c62_s_fa8), .Co(stage1_c62_c_fa8));
    FA fa_555(.A(stage0_r49_c13), .B(stage0_r50_c12), .C(stage0_r51_c11), .So(stage1_c62_s_fa9), .Co(stage1_c62_c_fa9));
    FA fa_556(.A(stage0_r52_c10), .B(stage0_r53_c9), .C(stage0_r54_c8), .So(stage1_c62_s_fa10), .Co(stage1_c62_c_fa10));
    FA fa_557(.A(stage0_r55_c7), .B(stage0_r56_c6), .C(stage0_r57_c5), .So(stage1_c62_s_fa11), .Co(stage1_c62_c_fa11));
    FA fa_558(.A(stage0_r58_c4), .B(stage0_r59_c3), .C(stage0_r60_c2), .So(stage1_c62_s_fa12), .Co(stage1_c62_c_fa12));
    HA ha_35(.A(stage0_r61_c1), .B(stage0_r62_c0), .So(stage1_c62_s_ha0), .Co(stage1_c62_c_ha0));
    FA fa_559(.A(stage0_r23_c40), .B(stage0_r24_c39), .C(stage0_r25_c38), .So(stage1_c63_s_fa0), .Co(stage1_c63_c_fa0));
    FA fa_560(.A(stage0_r26_c37), .B(stage0_r27_c36), .C(stage0_r28_c35), .So(stage1_c63_s_fa1), .Co(stage1_c63_c_fa1));
    FA fa_561(.A(stage0_r29_c34), .B(stage0_r30_c33), .C(stage0_r31_c32), .So(stage1_c63_s_fa2), .Co(stage1_c63_c_fa2));
    FA fa_562(.A(stage0_r32_c31), .B(stage0_r33_c30), .C(stage0_r34_c29), .So(stage1_c63_s_fa3), .Co(stage1_c63_c_fa3));
    FA fa_563(.A(stage0_r35_c28), .B(stage0_r36_c27), .C(stage0_r37_c26), .So(stage1_c63_s_fa4), .Co(stage1_c63_c_fa4));
    FA fa_564(.A(stage0_r38_c25), .B(stage0_r39_c24), .C(stage0_r40_c23), .So(stage1_c63_s_fa5), .Co(stage1_c63_c_fa5));
    FA fa_565(.A(stage0_r41_c22), .B(stage0_r42_c21), .C(stage0_r43_c20), .So(stage1_c63_s_fa6), .Co(stage1_c63_c_fa6));
    FA fa_566(.A(stage0_r44_c19), .B(stage0_r45_c18), .C(stage0_r46_c17), .So(stage1_c63_s_fa7), .Co(stage1_c63_c_fa7));
    FA fa_567(.A(stage0_r47_c16), .B(stage0_r48_c15), .C(stage0_r49_c14), .So(stage1_c63_s_fa8), .Co(stage1_c63_c_fa8));
    FA fa_568(.A(stage0_r50_c13), .B(stage0_r51_c12), .C(stage0_r52_c11), .So(stage1_c63_s_fa9), .Co(stage1_c63_c_fa9));
    FA fa_569(.A(stage0_r53_c10), .B(stage0_r54_c9), .C(stage0_r55_c8), .So(stage1_c63_s_fa10), .Co(stage1_c63_c_fa10));
    FA fa_570(.A(stage0_r56_c7), .B(stage0_r57_c6), .C(stage0_r58_c5), .So(stage1_c63_s_fa11), .Co(stage1_c63_c_fa11));
    FA fa_571(.A(stage0_r59_c4), .B(stage0_r60_c3), .C(stage0_r61_c2), .So(stage1_c63_s_fa12), .Co(stage1_c63_c_fa12));
    HA ha_36(.A(stage0_r62_c1), .B(stage0_r63_c0), .So(stage1_c63_s_ha0), .Co(stage1_c63_c_ha0));
    FA fa_572(.A(stage0_r24_c40), .B(stage0_r25_c39), .C(stage0_r26_c38), .So(stage1_c64_s_fa0), .Co(stage1_c64_c_fa0));
    FA fa_573(.A(stage0_r27_c37), .B(stage0_r28_c36), .C(stage0_r29_c35), .So(stage1_c64_s_fa1), .Co(stage1_c64_c_fa1));
    FA fa_574(.A(stage0_r30_c34), .B(stage0_r31_c33), .C(stage0_r32_c32), .So(stage1_c64_s_fa2), .Co(stage1_c64_c_fa2));
    FA fa_575(.A(stage0_r33_c31), .B(stage0_r34_c30), .C(stage0_r35_c29), .So(stage1_c64_s_fa3), .Co(stage1_c64_c_fa3));
    FA fa_576(.A(stage0_r36_c28), .B(stage0_r37_c27), .C(stage0_r38_c26), .So(stage1_c64_s_fa4), .Co(stage1_c64_c_fa4));
    FA fa_577(.A(stage0_r39_c25), .B(stage0_r40_c24), .C(stage0_r41_c23), .So(stage1_c64_s_fa5), .Co(stage1_c64_c_fa5));
    FA fa_578(.A(stage0_r42_c22), .B(stage0_r43_c21), .C(stage0_r44_c20), .So(stage1_c64_s_fa6), .Co(stage1_c64_c_fa6));
    FA fa_579(.A(stage0_r45_c19), .B(stage0_r46_c18), .C(stage0_r47_c17), .So(stage1_c64_s_fa7), .Co(stage1_c64_c_fa7));
    FA fa_580(.A(stage0_r48_c16), .B(stage0_r49_c15), .C(stage0_r50_c14), .So(stage1_c64_s_fa8), .Co(stage1_c64_c_fa8));
    FA fa_581(.A(stage0_r51_c13), .B(stage0_r52_c12), .C(stage0_r53_c11), .So(stage1_c64_s_fa9), .Co(stage1_c64_c_fa9));
    FA fa_582(.A(stage0_r54_c10), .B(stage0_r55_c9), .C(stage0_r56_c8), .So(stage1_c64_s_fa10), .Co(stage1_c64_c_fa10));
    FA fa_583(.A(stage0_r57_c7), .B(stage0_r58_c6), .C(stage0_r59_c5), .So(stage1_c64_s_fa11), .Co(stage1_c64_c_fa11));
    FA fa_584(.A(stage0_r60_c4), .B(stage0_r61_c3), .C(stage0_r62_c2), .So(stage1_c64_s_fa12), .Co(stage1_c64_c_fa12));
    HA ha_37(.A(stage0_r63_c1), .B(stage0_r64_c0), .So(stage1_c64_s_ha0), .Co(stage1_c64_c_ha0));
    FA fa_585(.A(stage0_r25_c40), .B(stage0_r26_c39), .C(stage0_r27_c38), .So(stage1_c65_s_fa0), .Co(stage1_c65_c_fa0));
    FA fa_586(.A(stage0_r28_c37), .B(stage0_r29_c36), .C(stage0_r30_c35), .So(stage1_c65_s_fa1), .Co(stage1_c65_c_fa1));
    FA fa_587(.A(stage0_r31_c34), .B(stage0_r32_c33), .C(stage0_r33_c32), .So(stage1_c65_s_fa2), .Co(stage1_c65_c_fa2));
    FA fa_588(.A(stage0_r34_c31), .B(stage0_r35_c30), .C(stage0_r36_c29), .So(stage1_c65_s_fa3), .Co(stage1_c65_c_fa3));
    FA fa_589(.A(stage0_r37_c28), .B(stage0_r38_c27), .C(stage0_r39_c26), .So(stage1_c65_s_fa4), .Co(stage1_c65_c_fa4));
    FA fa_590(.A(stage0_r40_c25), .B(stage0_r41_c24), .C(stage0_r42_c23), .So(stage1_c65_s_fa5), .Co(stage1_c65_c_fa5));
    FA fa_591(.A(stage0_r43_c22), .B(stage0_r44_c21), .C(stage0_r45_c20), .So(stage1_c65_s_fa6), .Co(stage1_c65_c_fa6));
    FA fa_592(.A(stage0_r46_c19), .B(stage0_r47_c18), .C(stage0_r48_c17), .So(stage1_c65_s_fa7), .Co(stage1_c65_c_fa7));
    FA fa_593(.A(stage0_r49_c16), .B(stage0_r50_c15), .C(stage0_r51_c14), .So(stage1_c65_s_fa8), .Co(stage1_c65_c_fa8));
    FA fa_594(.A(stage0_r52_c13), .B(stage0_r53_c12), .C(stage0_r54_c11), .So(stage1_c65_s_fa9), .Co(stage1_c65_c_fa9));
    FA fa_595(.A(stage0_r55_c10), .B(stage0_r56_c9), .C(stage0_r57_c8), .So(stage1_c65_s_fa10), .Co(stage1_c65_c_fa10));
    FA fa_596(.A(stage0_r58_c7), .B(stage0_r59_c6), .C(stage0_r60_c5), .So(stage1_c65_s_fa11), .Co(stage1_c65_c_fa11));
    FA fa_597(.A(stage0_r61_c4), .B(stage0_r62_c3), .C(stage0_r63_c2), .So(stage1_c65_s_fa12), .Co(stage1_c65_c_fa12));
    HA ha_38(.A(stage0_r64_c1), .B(stage0_r65_c0), .So(stage1_c65_s_ha0), .Co(stage1_c65_c_ha0));
    FA fa_598(.A(stage0_r26_c40), .B(stage0_r27_c39), .C(stage0_r28_c38), .So(stage1_c66_s_fa0), .Co(stage1_c66_c_fa0));
    FA fa_599(.A(stage0_r29_c37), .B(stage0_r30_c36), .C(stage0_r31_c35), .So(stage1_c66_s_fa1), .Co(stage1_c66_c_fa1));
    FA fa_600(.A(stage0_r32_c34), .B(stage0_r33_c33), .C(stage0_r34_c32), .So(stage1_c66_s_fa2), .Co(stage1_c66_c_fa2));
    FA fa_601(.A(stage0_r35_c31), .B(stage0_r36_c30), .C(stage0_r37_c29), .So(stage1_c66_s_fa3), .Co(stage1_c66_c_fa3));
    FA fa_602(.A(stage0_r38_c28), .B(stage0_r39_c27), .C(stage0_r40_c26), .So(stage1_c66_s_fa4), .Co(stage1_c66_c_fa4));
    FA fa_603(.A(stage0_r41_c25), .B(stage0_r42_c24), .C(stage0_r43_c23), .So(stage1_c66_s_fa5), .Co(stage1_c66_c_fa5));
    FA fa_604(.A(stage0_r44_c22), .B(stage0_r45_c21), .C(stage0_r46_c20), .So(stage1_c66_s_fa6), .Co(stage1_c66_c_fa6));
    FA fa_605(.A(stage0_r47_c19), .B(stage0_r48_c18), .C(stage0_r49_c17), .So(stage1_c66_s_fa7), .Co(stage1_c66_c_fa7));
    FA fa_606(.A(stage0_r50_c16), .B(stage0_r51_c15), .C(stage0_r52_c14), .So(stage1_c66_s_fa8), .Co(stage1_c66_c_fa8));
    FA fa_607(.A(stage0_r53_c13), .B(stage0_r54_c12), .C(stage0_r55_c11), .So(stage1_c66_s_fa9), .Co(stage1_c66_c_fa9));
    FA fa_608(.A(stage0_r56_c10), .B(stage0_r57_c9), .C(stage0_r58_c8), .So(stage1_c66_s_fa10), .Co(stage1_c66_c_fa10));
    FA fa_609(.A(stage0_r59_c7), .B(stage0_r60_c6), .C(stage0_r61_c5), .So(stage1_c66_s_fa11), .Co(stage1_c66_c_fa11));
    FA fa_610(.A(stage0_r62_c4), .B(stage0_r63_c3), .C(stage0_r64_c2), .So(stage1_c66_s_fa12), .Co(stage1_c66_c_fa12));
    HA ha_39(.A(stage0_r65_c1), .B(stage0_r66_c0), .So(stage1_c66_s_ha0), .Co(stage1_c66_c_ha0));
    FA fa_611(.A(stage0_r27_c40), .B(stage0_r28_c39), .C(stage0_r29_c38), .So(stage1_c67_s_fa0), .Co(stage1_c67_c_fa0));
    FA fa_612(.A(stage0_r30_c37), .B(stage0_r31_c36), .C(stage0_r32_c35), .So(stage1_c67_s_fa1), .Co(stage1_c67_c_fa1));
    FA fa_613(.A(stage0_r33_c34), .B(stage0_r34_c33), .C(stage0_r35_c32), .So(stage1_c67_s_fa2), .Co(stage1_c67_c_fa2));
    FA fa_614(.A(stage0_r36_c31), .B(stage0_r37_c30), .C(stage0_r38_c29), .So(stage1_c67_s_fa3), .Co(stage1_c67_c_fa3));
    FA fa_615(.A(stage0_r39_c28), .B(stage0_r40_c27), .C(stage0_r41_c26), .So(stage1_c67_s_fa4), .Co(stage1_c67_c_fa4));
    FA fa_616(.A(stage0_r42_c25), .B(stage0_r43_c24), .C(stage0_r44_c23), .So(stage1_c67_s_fa5), .Co(stage1_c67_c_fa5));
    FA fa_617(.A(stage0_r45_c22), .B(stage0_r46_c21), .C(stage0_r47_c20), .So(stage1_c67_s_fa6), .Co(stage1_c67_c_fa6));
    FA fa_618(.A(stage0_r48_c19), .B(stage0_r49_c18), .C(stage0_r50_c17), .So(stage1_c67_s_fa7), .Co(stage1_c67_c_fa7));
    FA fa_619(.A(stage0_r51_c16), .B(stage0_r52_c15), .C(stage0_r53_c14), .So(stage1_c67_s_fa8), .Co(stage1_c67_c_fa8));
    FA fa_620(.A(stage0_r54_c13), .B(stage0_r55_c12), .C(stage0_r56_c11), .So(stage1_c67_s_fa9), .Co(stage1_c67_c_fa9));
    FA fa_621(.A(stage0_r57_c10), .B(stage0_r58_c9), .C(stage0_r59_c8), .So(stage1_c67_s_fa10), .Co(stage1_c67_c_fa10));
    FA fa_622(.A(stage0_r60_c7), .B(stage0_r61_c6), .C(stage0_r62_c5), .So(stage1_c67_s_fa11), .Co(stage1_c67_c_fa11));
    FA fa_623(.A(stage0_r63_c4), .B(stage0_r64_c3), .C(stage0_r65_c2), .So(stage1_c67_s_fa12), .Co(stage1_c67_c_fa12));
    HA ha_40(.A(stage0_r66_c1), .B(stage0_r67_c0), .So(stage1_c67_s_ha0), .Co(stage1_c67_c_ha0));
    FA fa_624(.A(stage0_r28_c40), .B(stage0_r29_c39), .C(stage0_r30_c38), .So(stage1_c68_s_fa0), .Co(stage1_c68_c_fa0));
    FA fa_625(.A(stage0_r31_c37), .B(stage0_r32_c36), .C(stage0_r33_c35), .So(stage1_c68_s_fa1), .Co(stage1_c68_c_fa1));
    FA fa_626(.A(stage0_r34_c34), .B(stage0_r35_c33), .C(stage0_r36_c32), .So(stage1_c68_s_fa2), .Co(stage1_c68_c_fa2));
    FA fa_627(.A(stage0_r37_c31), .B(stage0_r38_c30), .C(stage0_r39_c29), .So(stage1_c68_s_fa3), .Co(stage1_c68_c_fa3));
    FA fa_628(.A(stage0_r40_c28), .B(stage0_r41_c27), .C(stage0_r42_c26), .So(stage1_c68_s_fa4), .Co(stage1_c68_c_fa4));
    FA fa_629(.A(stage0_r43_c25), .B(stage0_r44_c24), .C(stage0_r45_c23), .So(stage1_c68_s_fa5), .Co(stage1_c68_c_fa5));
    FA fa_630(.A(stage0_r46_c22), .B(stage0_r47_c21), .C(stage0_r48_c20), .So(stage1_c68_s_fa6), .Co(stage1_c68_c_fa6));
    FA fa_631(.A(stage0_r49_c19), .B(stage0_r50_c18), .C(stage0_r51_c17), .So(stage1_c68_s_fa7), .Co(stage1_c68_c_fa7));
    FA fa_632(.A(stage0_r52_c16), .B(stage0_r53_c15), .C(stage0_r54_c14), .So(stage1_c68_s_fa8), .Co(stage1_c68_c_fa8));
    FA fa_633(.A(stage0_r55_c13), .B(stage0_r56_c12), .C(stage0_r57_c11), .So(stage1_c68_s_fa9), .Co(stage1_c68_c_fa9));
    FA fa_634(.A(stage0_r58_c10), .B(stage0_r59_c9), .C(stage0_r60_c8), .So(stage1_c68_s_fa10), .Co(stage1_c68_c_fa10));
    FA fa_635(.A(stage0_r61_c7), .B(stage0_r62_c6), .C(stage0_r63_c5), .So(stage1_c68_s_fa11), .Co(stage1_c68_c_fa11));
    FA fa_636(.A(stage0_r64_c4), .B(stage0_r65_c3), .C(stage0_r66_c2), .So(stage1_c68_s_fa12), .Co(stage1_c68_c_fa12));
    HA ha_41(.A(stage0_r67_c1), .B(stage0_r68_c0), .So(stage1_c68_s_ha0), .Co(stage1_c68_c_ha0));
    FA fa_637(.A(stage0_r29_c40), .B(stage0_r30_c39), .C(stage0_r31_c38), .So(stage1_c69_s_fa0), .Co(stage1_c69_c_fa0));
    FA fa_638(.A(stage0_r32_c37), .B(stage0_r33_c36), .C(stage0_r34_c35), .So(stage1_c69_s_fa1), .Co(stage1_c69_c_fa1));
    FA fa_639(.A(stage0_r35_c34), .B(stage0_r36_c33), .C(stage0_r37_c32), .So(stage1_c69_s_fa2), .Co(stage1_c69_c_fa2));
    FA fa_640(.A(stage0_r38_c31), .B(stage0_r39_c30), .C(stage0_r40_c29), .So(stage1_c69_s_fa3), .Co(stage1_c69_c_fa3));
    FA fa_641(.A(stage0_r41_c28), .B(stage0_r42_c27), .C(stage0_r43_c26), .So(stage1_c69_s_fa4), .Co(stage1_c69_c_fa4));
    FA fa_642(.A(stage0_r44_c25), .B(stage0_r45_c24), .C(stage0_r46_c23), .So(stage1_c69_s_fa5), .Co(stage1_c69_c_fa5));
    FA fa_643(.A(stage0_r47_c22), .B(stage0_r48_c21), .C(stage0_r49_c20), .So(stage1_c69_s_fa6), .Co(stage1_c69_c_fa6));
    FA fa_644(.A(stage0_r50_c19), .B(stage0_r51_c18), .C(stage0_r52_c17), .So(stage1_c69_s_fa7), .Co(stage1_c69_c_fa7));
    FA fa_645(.A(stage0_r53_c16), .B(stage0_r54_c15), .C(stage0_r55_c14), .So(stage1_c69_s_fa8), .Co(stage1_c69_c_fa8));
    FA fa_646(.A(stage0_r56_c13), .B(stage0_r57_c12), .C(stage0_r58_c11), .So(stage1_c69_s_fa9), .Co(stage1_c69_c_fa9));
    FA fa_647(.A(stage0_r59_c10), .B(stage0_r60_c9), .C(stage0_r61_c8), .So(stage1_c69_s_fa10), .Co(stage1_c69_c_fa10));
    FA fa_648(.A(stage0_r62_c7), .B(stage0_r63_c6), .C(stage0_r64_c5), .So(stage1_c69_s_fa11), .Co(stage1_c69_c_fa11));
    FA fa_649(.A(stage0_r65_c4), .B(stage0_r66_c3), .C(stage0_r67_c2), .So(stage1_c69_s_fa12), .Co(stage1_c69_c_fa12));
    HA ha_42(.A(stage0_r68_c1), .B(stage0_r69_c0), .So(stage1_c69_s_ha0), .Co(stage1_c69_c_ha0));
    FA fa_650(.A(stage0_r30_c40), .B(stage0_r31_c39), .C(stage0_r32_c38), .So(stage1_c70_s_fa0), .Co(stage1_c70_c_fa0));
    FA fa_651(.A(stage0_r33_c37), .B(stage0_r34_c36), .C(stage0_r35_c35), .So(stage1_c70_s_fa1), .Co(stage1_c70_c_fa1));
    FA fa_652(.A(stage0_r36_c34), .B(stage0_r37_c33), .C(stage0_r38_c32), .So(stage1_c70_s_fa2), .Co(stage1_c70_c_fa2));
    FA fa_653(.A(stage0_r39_c31), .B(stage0_r40_c30), .C(stage0_r41_c29), .So(stage1_c70_s_fa3), .Co(stage1_c70_c_fa3));
    FA fa_654(.A(stage0_r42_c28), .B(stage0_r43_c27), .C(stage0_r44_c26), .So(stage1_c70_s_fa4), .Co(stage1_c70_c_fa4));
    FA fa_655(.A(stage0_r45_c25), .B(stage0_r46_c24), .C(stage0_r47_c23), .So(stage1_c70_s_fa5), .Co(stage1_c70_c_fa5));
    FA fa_656(.A(stage0_r48_c22), .B(stage0_r49_c21), .C(stage0_r50_c20), .So(stage1_c70_s_fa6), .Co(stage1_c70_c_fa6));
    FA fa_657(.A(stage0_r51_c19), .B(stage0_r52_c18), .C(stage0_r53_c17), .So(stage1_c70_s_fa7), .Co(stage1_c70_c_fa7));
    FA fa_658(.A(stage0_r54_c16), .B(stage0_r55_c15), .C(stage0_r56_c14), .So(stage1_c70_s_fa8), .Co(stage1_c70_c_fa8));
    FA fa_659(.A(stage0_r57_c13), .B(stage0_r58_c12), .C(stage0_r59_c11), .So(stage1_c70_s_fa9), .Co(stage1_c70_c_fa9));
    FA fa_660(.A(stage0_r60_c10), .B(stage0_r61_c9), .C(stage0_r62_c8), .So(stage1_c70_s_fa10), .Co(stage1_c70_c_fa10));
    FA fa_661(.A(stage0_r63_c7), .B(stage0_r64_c6), .C(stage0_r65_c5), .So(stage1_c70_s_fa11), .Co(stage1_c70_c_fa11));
    FA fa_662(.A(stage0_r66_c4), .B(stage0_r67_c3), .C(stage0_r68_c2), .So(stage1_c70_s_fa12), .Co(stage1_c70_c_fa12));
    HA ha_43(.A(stage0_r69_c1), .B(stage0_r70_c0), .So(stage1_c70_s_ha0), .Co(stage1_c70_c_ha0));
    FA fa_663(.A(stage0_r31_c40), .B(stage0_r32_c39), .C(stage0_r33_c38), .So(stage1_c71_s_fa0), .Co(stage1_c71_c_fa0));
    FA fa_664(.A(stage0_r34_c37), .B(stage0_r35_c36), .C(stage0_r36_c35), .So(stage1_c71_s_fa1), .Co(stage1_c71_c_fa1));
    FA fa_665(.A(stage0_r37_c34), .B(stage0_r38_c33), .C(stage0_r39_c32), .So(stage1_c71_s_fa2), .Co(stage1_c71_c_fa2));
    FA fa_666(.A(stage0_r40_c31), .B(stage0_r41_c30), .C(stage0_r42_c29), .So(stage1_c71_s_fa3), .Co(stage1_c71_c_fa3));
    FA fa_667(.A(stage0_r43_c28), .B(stage0_r44_c27), .C(stage0_r45_c26), .So(stage1_c71_s_fa4), .Co(stage1_c71_c_fa4));
    FA fa_668(.A(stage0_r46_c25), .B(stage0_r47_c24), .C(stage0_r48_c23), .So(stage1_c71_s_fa5), .Co(stage1_c71_c_fa5));
    FA fa_669(.A(stage0_r49_c22), .B(stage0_r50_c21), .C(stage0_r51_c20), .So(stage1_c71_s_fa6), .Co(stage1_c71_c_fa6));
    FA fa_670(.A(stage0_r52_c19), .B(stage0_r53_c18), .C(stage0_r54_c17), .So(stage1_c71_s_fa7), .Co(stage1_c71_c_fa7));
    FA fa_671(.A(stage0_r55_c16), .B(stage0_r56_c15), .C(stage0_r57_c14), .So(stage1_c71_s_fa8), .Co(stage1_c71_c_fa8));
    FA fa_672(.A(stage0_r58_c13), .B(stage0_r59_c12), .C(stage0_r60_c11), .So(stage1_c71_s_fa9), .Co(stage1_c71_c_fa9));
    FA fa_673(.A(stage0_r61_c10), .B(stage0_r62_c9), .C(stage0_r63_c8), .So(stage1_c71_s_fa10), .Co(stage1_c71_c_fa10));
    FA fa_674(.A(stage0_r64_c7), .B(stage0_r65_c6), .C(stage0_r66_c5), .So(stage1_c71_s_fa11), .Co(stage1_c71_c_fa11));
    FA fa_675(.A(stage0_r67_c4), .B(stage0_r68_c3), .C(stage0_r69_c2), .So(stage1_c71_s_fa12), .Co(stage1_c71_c_fa12));
    HA ha_44(.A(stage0_r70_c1), .B(stage0_r71_c0), .So(stage1_c71_s_ha0), .Co(stage1_c71_c_ha0));
    FA fa_676(.A(stage0_r32_c40), .B(stage0_r33_c39), .C(stage0_r34_c38), .So(stage1_c72_s_fa0), .Co(stage1_c72_c_fa0));
    FA fa_677(.A(stage0_r35_c37), .B(stage0_r36_c36), .C(stage0_r37_c35), .So(stage1_c72_s_fa1), .Co(stage1_c72_c_fa1));
    FA fa_678(.A(stage0_r38_c34), .B(stage0_r39_c33), .C(stage0_r40_c32), .So(stage1_c72_s_fa2), .Co(stage1_c72_c_fa2));
    FA fa_679(.A(stage0_r41_c31), .B(stage0_r42_c30), .C(stage0_r43_c29), .So(stage1_c72_s_fa3), .Co(stage1_c72_c_fa3));
    FA fa_680(.A(stage0_r44_c28), .B(stage0_r45_c27), .C(stage0_r46_c26), .So(stage1_c72_s_fa4), .Co(stage1_c72_c_fa4));
    FA fa_681(.A(stage0_r47_c25), .B(stage0_r48_c24), .C(stage0_r49_c23), .So(stage1_c72_s_fa5), .Co(stage1_c72_c_fa5));
    FA fa_682(.A(stage0_r50_c22), .B(stage0_r51_c21), .C(stage0_r52_c20), .So(stage1_c72_s_fa6), .Co(stage1_c72_c_fa6));
    FA fa_683(.A(stage0_r53_c19), .B(stage0_r54_c18), .C(stage0_r55_c17), .So(stage1_c72_s_fa7), .Co(stage1_c72_c_fa7));
    FA fa_684(.A(stage0_r56_c16), .B(stage0_r57_c15), .C(stage0_r58_c14), .So(stage1_c72_s_fa8), .Co(stage1_c72_c_fa8));
    FA fa_685(.A(stage0_r59_c13), .B(stage0_r60_c12), .C(stage0_r61_c11), .So(stage1_c72_s_fa9), .Co(stage1_c72_c_fa9));
    FA fa_686(.A(stage0_r62_c10), .B(stage0_r63_c9), .C(stage0_r64_c8), .So(stage1_c72_s_fa10), .Co(stage1_c72_c_fa10));
    FA fa_687(.A(stage0_r65_c7), .B(stage0_r66_c6), .C(stage0_r67_c5), .So(stage1_c72_s_fa11), .Co(stage1_c72_c_fa11));
    FA fa_688(.A(stage0_r68_c4), .B(stage0_r69_c3), .C(stage0_r70_c2), .So(stage1_c72_s_fa12), .Co(stage1_c72_c_fa12));
    FA fa_689(.A(stage0_r33_c40), .B(stage0_r34_c39), .C(stage0_r35_c38), .So(stage1_c73_s_fa0), .Co(stage1_c73_c_fa0));
    FA fa_690(.A(stage0_r36_c37), .B(stage0_r37_c36), .C(stage0_r38_c35), .So(stage1_c73_s_fa1), .Co(stage1_c73_c_fa1));
    FA fa_691(.A(stage0_r39_c34), .B(stage0_r40_c33), .C(stage0_r41_c32), .So(stage1_c73_s_fa2), .Co(stage1_c73_c_fa2));
    FA fa_692(.A(stage0_r42_c31), .B(stage0_r43_c30), .C(stage0_r44_c29), .So(stage1_c73_s_fa3), .Co(stage1_c73_c_fa3));
    FA fa_693(.A(stage0_r45_c28), .B(stage0_r46_c27), .C(stage0_r47_c26), .So(stage1_c73_s_fa4), .Co(stage1_c73_c_fa4));
    FA fa_694(.A(stage0_r48_c25), .B(stage0_r49_c24), .C(stage0_r50_c23), .So(stage1_c73_s_fa5), .Co(stage1_c73_c_fa5));
    FA fa_695(.A(stage0_r51_c22), .B(stage0_r52_c21), .C(stage0_r53_c20), .So(stage1_c73_s_fa6), .Co(stage1_c73_c_fa6));
    FA fa_696(.A(stage0_r54_c19), .B(stage0_r55_c18), .C(stage0_r56_c17), .So(stage1_c73_s_fa7), .Co(stage1_c73_c_fa7));
    FA fa_697(.A(stage0_r57_c16), .B(stage0_r58_c15), .C(stage0_r59_c14), .So(stage1_c73_s_fa8), .Co(stage1_c73_c_fa8));
    FA fa_698(.A(stage0_r60_c13), .B(stage0_r61_c12), .C(stage0_r62_c11), .So(stage1_c73_s_fa9), .Co(stage1_c73_c_fa9));
    FA fa_699(.A(stage0_r63_c10), .B(stage0_r64_c9), .C(stage0_r65_c8), .So(stage1_c73_s_fa10), .Co(stage1_c73_c_fa10));
    FA fa_700(.A(stage0_r66_c7), .B(stage0_r67_c6), .C(stage0_r68_c5), .So(stage1_c73_s_fa11), .Co(stage1_c73_c_fa11));
    FA fa_701(.A(stage0_r69_c4), .B(stage0_r70_c3), .C(stage0_r71_c2), .So(stage1_c73_s_fa12), .Co(stage1_c73_c_fa12));
    FA fa_702(.A(stage0_r34_c40), .B(stage0_r35_c39), .C(stage0_r36_c38), .So(stage1_c74_s_fa0), .Co(stage1_c74_c_fa0));
    FA fa_703(.A(stage0_r37_c37), .B(stage0_r38_c36), .C(stage0_r39_c35), .So(stage1_c74_s_fa1), .Co(stage1_c74_c_fa1));
    FA fa_704(.A(stage0_r40_c34), .B(stage0_r41_c33), .C(stage0_r42_c32), .So(stage1_c74_s_fa2), .Co(stage1_c74_c_fa2));
    FA fa_705(.A(stage0_r43_c31), .B(stage0_r44_c30), .C(stage0_r45_c29), .So(stage1_c74_s_fa3), .Co(stage1_c74_c_fa3));
    FA fa_706(.A(stage0_r46_c28), .B(stage0_r47_c27), .C(stage0_r48_c26), .So(stage1_c74_s_fa4), .Co(stage1_c74_c_fa4));
    FA fa_707(.A(stage0_r49_c25), .B(stage0_r50_c24), .C(stage0_r51_c23), .So(stage1_c74_s_fa5), .Co(stage1_c74_c_fa5));
    FA fa_708(.A(stage0_r52_c22), .B(stage0_r53_c21), .C(stage0_r54_c20), .So(stage1_c74_s_fa6), .Co(stage1_c74_c_fa6));
    FA fa_709(.A(stage0_r55_c19), .B(stage0_r56_c18), .C(stage0_r57_c17), .So(stage1_c74_s_fa7), .Co(stage1_c74_c_fa7));
    FA fa_710(.A(stage0_r58_c16), .B(stage0_r59_c15), .C(stage0_r60_c14), .So(stage1_c74_s_fa8), .Co(stage1_c74_c_fa8));
    FA fa_711(.A(stage0_r61_c13), .B(stage0_r62_c12), .C(stage0_r63_c11), .So(stage1_c74_s_fa9), .Co(stage1_c74_c_fa9));
    FA fa_712(.A(stage0_r64_c10), .B(stage0_r65_c9), .C(stage0_r66_c8), .So(stage1_c74_s_fa10), .Co(stage1_c74_c_fa10));
    FA fa_713(.A(stage0_r67_c7), .B(stage0_r68_c6), .C(stage0_r69_c5), .So(stage1_c74_s_fa11), .Co(stage1_c74_c_fa11));
    HA ha_45(.A(stage0_r70_c4), .B(stage0_r71_c3), .So(stage1_c74_s_ha0), .Co(stage1_c74_c_ha0));
    FA fa_714(.A(stage0_r35_c40), .B(stage0_r36_c39), .C(stage0_r37_c38), .So(stage1_c75_s_fa0), .Co(stage1_c75_c_fa0));
    FA fa_715(.A(stage0_r38_c37), .B(stage0_r39_c36), .C(stage0_r40_c35), .So(stage1_c75_s_fa1), .Co(stage1_c75_c_fa1));
    FA fa_716(.A(stage0_r41_c34), .B(stage0_r42_c33), .C(stage0_r43_c32), .So(stage1_c75_s_fa2), .Co(stage1_c75_c_fa2));
    FA fa_717(.A(stage0_r44_c31), .B(stage0_r45_c30), .C(stage0_r46_c29), .So(stage1_c75_s_fa3), .Co(stage1_c75_c_fa3));
    FA fa_718(.A(stage0_r47_c28), .B(stage0_r48_c27), .C(stage0_r49_c26), .So(stage1_c75_s_fa4), .Co(stage1_c75_c_fa4));
    FA fa_719(.A(stage0_r50_c25), .B(stage0_r51_c24), .C(stage0_r52_c23), .So(stage1_c75_s_fa5), .Co(stage1_c75_c_fa5));
    FA fa_720(.A(stage0_r53_c22), .B(stage0_r54_c21), .C(stage0_r55_c20), .So(stage1_c75_s_fa6), .Co(stage1_c75_c_fa6));
    FA fa_721(.A(stage0_r56_c19), .B(stage0_r57_c18), .C(stage0_r58_c17), .So(stage1_c75_s_fa7), .Co(stage1_c75_c_fa7));
    FA fa_722(.A(stage0_r59_c16), .B(stage0_r60_c15), .C(stage0_r61_c14), .So(stage1_c75_s_fa8), .Co(stage1_c75_c_fa8));
    FA fa_723(.A(stage0_r62_c13), .B(stage0_r63_c12), .C(stage0_r64_c11), .So(stage1_c75_s_fa9), .Co(stage1_c75_c_fa9));
    FA fa_724(.A(stage0_r65_c10), .B(stage0_r66_c9), .C(stage0_r67_c8), .So(stage1_c75_s_fa10), .Co(stage1_c75_c_fa10));
    FA fa_725(.A(stage0_r68_c7), .B(stage0_r69_c6), .C(stage0_r70_c5), .So(stage1_c75_s_fa11), .Co(stage1_c75_c_fa11));
    FA fa_726(.A(stage0_r36_c40), .B(stage0_r37_c39), .C(stage0_r38_c38), .So(stage1_c76_s_fa0), .Co(stage1_c76_c_fa0));
    FA fa_727(.A(stage0_r39_c37), .B(stage0_r40_c36), .C(stage0_r41_c35), .So(stage1_c76_s_fa1), .Co(stage1_c76_c_fa1));
    FA fa_728(.A(stage0_r42_c34), .B(stage0_r43_c33), .C(stage0_r44_c32), .So(stage1_c76_s_fa2), .Co(stage1_c76_c_fa2));
    FA fa_729(.A(stage0_r45_c31), .B(stage0_r46_c30), .C(stage0_r47_c29), .So(stage1_c76_s_fa3), .Co(stage1_c76_c_fa3));
    FA fa_730(.A(stage0_r48_c28), .B(stage0_r49_c27), .C(stage0_r50_c26), .So(stage1_c76_s_fa4), .Co(stage1_c76_c_fa4));
    FA fa_731(.A(stage0_r51_c25), .B(stage0_r52_c24), .C(stage0_r53_c23), .So(stage1_c76_s_fa5), .Co(stage1_c76_c_fa5));
    FA fa_732(.A(stage0_r54_c22), .B(stage0_r55_c21), .C(stage0_r56_c20), .So(stage1_c76_s_fa6), .Co(stage1_c76_c_fa6));
    FA fa_733(.A(stage0_r57_c19), .B(stage0_r58_c18), .C(stage0_r59_c17), .So(stage1_c76_s_fa7), .Co(stage1_c76_c_fa7));
    FA fa_734(.A(stage0_r60_c16), .B(stage0_r61_c15), .C(stage0_r62_c14), .So(stage1_c76_s_fa8), .Co(stage1_c76_c_fa8));
    FA fa_735(.A(stage0_r63_c13), .B(stage0_r64_c12), .C(stage0_r65_c11), .So(stage1_c76_s_fa9), .Co(stage1_c76_c_fa9));
    FA fa_736(.A(stage0_r66_c10), .B(stage0_r67_c9), .C(stage0_r68_c8), .So(stage1_c76_s_fa10), .Co(stage1_c76_c_fa10));
    FA fa_737(.A(stage0_r69_c7), .B(stage0_r70_c6), .C(stage0_r71_c5), .So(stage1_c76_s_fa11), .Co(stage1_c76_c_fa11));
    FA fa_738(.A(stage0_r37_c40), .B(stage0_r38_c39), .C(stage0_r39_c38), .So(stage1_c77_s_fa0), .Co(stage1_c77_c_fa0));
    FA fa_739(.A(stage0_r40_c37), .B(stage0_r41_c36), .C(stage0_r42_c35), .So(stage1_c77_s_fa1), .Co(stage1_c77_c_fa1));
    FA fa_740(.A(stage0_r43_c34), .B(stage0_r44_c33), .C(stage0_r45_c32), .So(stage1_c77_s_fa2), .Co(stage1_c77_c_fa2));
    FA fa_741(.A(stage0_r46_c31), .B(stage0_r47_c30), .C(stage0_r48_c29), .So(stage1_c77_s_fa3), .Co(stage1_c77_c_fa3));
    FA fa_742(.A(stage0_r49_c28), .B(stage0_r50_c27), .C(stage0_r51_c26), .So(stage1_c77_s_fa4), .Co(stage1_c77_c_fa4));
    FA fa_743(.A(stage0_r52_c25), .B(stage0_r53_c24), .C(stage0_r54_c23), .So(stage1_c77_s_fa5), .Co(stage1_c77_c_fa5));
    FA fa_744(.A(stage0_r55_c22), .B(stage0_r56_c21), .C(stage0_r57_c20), .So(stage1_c77_s_fa6), .Co(stage1_c77_c_fa6));
    FA fa_745(.A(stage0_r58_c19), .B(stage0_r59_c18), .C(stage0_r60_c17), .So(stage1_c77_s_fa7), .Co(stage1_c77_c_fa7));
    FA fa_746(.A(stage0_r61_c16), .B(stage0_r62_c15), .C(stage0_r63_c14), .So(stage1_c77_s_fa8), .Co(stage1_c77_c_fa8));
    FA fa_747(.A(stage0_r64_c13), .B(stage0_r65_c12), .C(stage0_r66_c11), .So(stage1_c77_s_fa9), .Co(stage1_c77_c_fa9));
    FA fa_748(.A(stage0_r67_c10), .B(stage0_r68_c9), .C(stage0_r69_c8), .So(stage1_c77_s_fa10), .Co(stage1_c77_c_fa10));
    HA ha_46(.A(stage0_r70_c7), .B(stage0_r71_c6), .So(stage1_c77_s_ha0), .Co(stage1_c77_c_ha0));
    FA fa_749(.A(stage0_r38_c40), .B(stage0_r39_c39), .C(stage0_r40_c38), .So(stage1_c78_s_fa0), .Co(stage1_c78_c_fa0));
    FA fa_750(.A(stage0_r41_c37), .B(stage0_r42_c36), .C(stage0_r43_c35), .So(stage1_c78_s_fa1), .Co(stage1_c78_c_fa1));
    FA fa_751(.A(stage0_r44_c34), .B(stage0_r45_c33), .C(stage0_r46_c32), .So(stage1_c78_s_fa2), .Co(stage1_c78_c_fa2));
    FA fa_752(.A(stage0_r47_c31), .B(stage0_r48_c30), .C(stage0_r49_c29), .So(stage1_c78_s_fa3), .Co(stage1_c78_c_fa3));
    FA fa_753(.A(stage0_r50_c28), .B(stage0_r51_c27), .C(stage0_r52_c26), .So(stage1_c78_s_fa4), .Co(stage1_c78_c_fa4));
    FA fa_754(.A(stage0_r53_c25), .B(stage0_r54_c24), .C(stage0_r55_c23), .So(stage1_c78_s_fa5), .Co(stage1_c78_c_fa5));
    FA fa_755(.A(stage0_r56_c22), .B(stage0_r57_c21), .C(stage0_r58_c20), .So(stage1_c78_s_fa6), .Co(stage1_c78_c_fa6));
    FA fa_756(.A(stage0_r59_c19), .B(stage0_r60_c18), .C(stage0_r61_c17), .So(stage1_c78_s_fa7), .Co(stage1_c78_c_fa7));
    FA fa_757(.A(stage0_r62_c16), .B(stage0_r63_c15), .C(stage0_r64_c14), .So(stage1_c78_s_fa8), .Co(stage1_c78_c_fa8));
    FA fa_758(.A(stage0_r65_c13), .B(stage0_r66_c12), .C(stage0_r67_c11), .So(stage1_c78_s_fa9), .Co(stage1_c78_c_fa9));
    FA fa_759(.A(stage0_r68_c10), .B(stage0_r69_c9), .C(stage0_r70_c8), .So(stage1_c78_s_fa10), .Co(stage1_c78_c_fa10));
    FA fa_760(.A(stage0_r39_c40), .B(stage0_r40_c39), .C(stage0_r41_c38), .So(stage1_c79_s_fa0), .Co(stage1_c79_c_fa0));
    FA fa_761(.A(stage0_r42_c37), .B(stage0_r43_c36), .C(stage0_r44_c35), .So(stage1_c79_s_fa1), .Co(stage1_c79_c_fa1));
    FA fa_762(.A(stage0_r45_c34), .B(stage0_r46_c33), .C(stage0_r47_c32), .So(stage1_c79_s_fa2), .Co(stage1_c79_c_fa2));
    FA fa_763(.A(stage0_r48_c31), .B(stage0_r49_c30), .C(stage0_r50_c29), .So(stage1_c79_s_fa3), .Co(stage1_c79_c_fa3));
    FA fa_764(.A(stage0_r51_c28), .B(stage0_r52_c27), .C(stage0_r53_c26), .So(stage1_c79_s_fa4), .Co(stage1_c79_c_fa4));
    FA fa_765(.A(stage0_r54_c25), .B(stage0_r55_c24), .C(stage0_r56_c23), .So(stage1_c79_s_fa5), .Co(stage1_c79_c_fa5));
    FA fa_766(.A(stage0_r57_c22), .B(stage0_r58_c21), .C(stage0_r59_c20), .So(stage1_c79_s_fa6), .Co(stage1_c79_c_fa6));
    FA fa_767(.A(stage0_r60_c19), .B(stage0_r61_c18), .C(stage0_r62_c17), .So(stage1_c79_s_fa7), .Co(stage1_c79_c_fa7));
    FA fa_768(.A(stage0_r63_c16), .B(stage0_r64_c15), .C(stage0_r65_c14), .So(stage1_c79_s_fa8), .Co(stage1_c79_c_fa8));
    FA fa_769(.A(stage0_r66_c13), .B(stage0_r67_c12), .C(stage0_r68_c11), .So(stage1_c79_s_fa9), .Co(stage1_c79_c_fa9));
    FA fa_770(.A(stage0_r69_c10), .B(stage0_r70_c9), .C(stage0_r71_c8), .So(stage1_c79_s_fa10), .Co(stage1_c79_c_fa10));
    FA fa_771(.A(stage0_r40_c40), .B(stage0_r41_c39), .C(stage0_r42_c38), .So(stage1_c80_s_fa0), .Co(stage1_c80_c_fa0));
    FA fa_772(.A(stage0_r43_c37), .B(stage0_r44_c36), .C(stage0_r45_c35), .So(stage1_c80_s_fa1), .Co(stage1_c80_c_fa1));
    FA fa_773(.A(stage0_r46_c34), .B(stage0_r47_c33), .C(stage0_r48_c32), .So(stage1_c80_s_fa2), .Co(stage1_c80_c_fa2));
    FA fa_774(.A(stage0_r49_c31), .B(stage0_r50_c30), .C(stage0_r51_c29), .So(stage1_c80_s_fa3), .Co(stage1_c80_c_fa3));
    FA fa_775(.A(stage0_r52_c28), .B(stage0_r53_c27), .C(stage0_r54_c26), .So(stage1_c80_s_fa4), .Co(stage1_c80_c_fa4));
    FA fa_776(.A(stage0_r55_c25), .B(stage0_r56_c24), .C(stage0_r57_c23), .So(stage1_c80_s_fa5), .Co(stage1_c80_c_fa5));
    FA fa_777(.A(stage0_r58_c22), .B(stage0_r59_c21), .C(stage0_r60_c20), .So(stage1_c80_s_fa6), .Co(stage1_c80_c_fa6));
    FA fa_778(.A(stage0_r61_c19), .B(stage0_r62_c18), .C(stage0_r63_c17), .So(stage1_c80_s_fa7), .Co(stage1_c80_c_fa7));
    FA fa_779(.A(stage0_r64_c16), .B(stage0_r65_c15), .C(stage0_r66_c14), .So(stage1_c80_s_fa8), .Co(stage1_c80_c_fa8));
    FA fa_780(.A(stage0_r67_c13), .B(stage0_r68_c12), .C(stage0_r69_c11), .So(stage1_c80_s_fa9), .Co(stage1_c80_c_fa9));
    HA ha_47(.A(stage0_r70_c10), .B(stage0_r71_c9), .So(stage1_c80_s_ha0), .Co(stage1_c80_c_ha0));
    FA fa_781(.A(stage0_r41_c40), .B(stage0_r42_c39), .C(stage0_r43_c38), .So(stage1_c81_s_fa0), .Co(stage1_c81_c_fa0));
    FA fa_782(.A(stage0_r44_c37), .B(stage0_r45_c36), .C(stage0_r46_c35), .So(stage1_c81_s_fa1), .Co(stage1_c81_c_fa1));
    FA fa_783(.A(stage0_r47_c34), .B(stage0_r48_c33), .C(stage0_r49_c32), .So(stage1_c81_s_fa2), .Co(stage1_c81_c_fa2));
    FA fa_784(.A(stage0_r50_c31), .B(stage0_r51_c30), .C(stage0_r52_c29), .So(stage1_c81_s_fa3), .Co(stage1_c81_c_fa3));
    FA fa_785(.A(stage0_r53_c28), .B(stage0_r54_c27), .C(stage0_r55_c26), .So(stage1_c81_s_fa4), .Co(stage1_c81_c_fa4));
    FA fa_786(.A(stage0_r56_c25), .B(stage0_r57_c24), .C(stage0_r58_c23), .So(stage1_c81_s_fa5), .Co(stage1_c81_c_fa5));
    FA fa_787(.A(stage0_r59_c22), .B(stage0_r60_c21), .C(stage0_r61_c20), .So(stage1_c81_s_fa6), .Co(stage1_c81_c_fa6));
    FA fa_788(.A(stage0_r62_c19), .B(stage0_r63_c18), .C(stage0_r64_c17), .So(stage1_c81_s_fa7), .Co(stage1_c81_c_fa7));
    FA fa_789(.A(stage0_r65_c16), .B(stage0_r66_c15), .C(stage0_r67_c14), .So(stage1_c81_s_fa8), .Co(stage1_c81_c_fa8));
    FA fa_790(.A(stage0_r68_c13), .B(stage0_r69_c12), .C(stage0_r70_c11), .So(stage1_c81_s_fa9), .Co(stage1_c81_c_fa9));
    FA fa_791(.A(stage0_r42_c40), .B(stage0_r43_c39), .C(stage0_r44_c38), .So(stage1_c82_s_fa0), .Co(stage1_c82_c_fa0));
    FA fa_792(.A(stage0_r45_c37), .B(stage0_r46_c36), .C(stage0_r47_c35), .So(stage1_c82_s_fa1), .Co(stage1_c82_c_fa1));
    FA fa_793(.A(stage0_r48_c34), .B(stage0_r49_c33), .C(stage0_r50_c32), .So(stage1_c82_s_fa2), .Co(stage1_c82_c_fa2));
    FA fa_794(.A(stage0_r51_c31), .B(stage0_r52_c30), .C(stage0_r53_c29), .So(stage1_c82_s_fa3), .Co(stage1_c82_c_fa3));
    FA fa_795(.A(stage0_r54_c28), .B(stage0_r55_c27), .C(stage0_r56_c26), .So(stage1_c82_s_fa4), .Co(stage1_c82_c_fa4));
    FA fa_796(.A(stage0_r57_c25), .B(stage0_r58_c24), .C(stage0_r59_c23), .So(stage1_c82_s_fa5), .Co(stage1_c82_c_fa5));
    FA fa_797(.A(stage0_r60_c22), .B(stage0_r61_c21), .C(stage0_r62_c20), .So(stage1_c82_s_fa6), .Co(stage1_c82_c_fa6));
    FA fa_798(.A(stage0_r63_c19), .B(stage0_r64_c18), .C(stage0_r65_c17), .So(stage1_c82_s_fa7), .Co(stage1_c82_c_fa7));
    FA fa_799(.A(stage0_r66_c16), .B(stage0_r67_c15), .C(stage0_r68_c14), .So(stage1_c82_s_fa8), .Co(stage1_c82_c_fa8));
    FA fa_800(.A(stage0_r69_c13), .B(stage0_r70_c12), .C(stage0_r71_c11), .So(stage1_c82_s_fa9), .Co(stage1_c82_c_fa9));
    FA fa_801(.A(stage0_r43_c40), .B(stage0_r44_c39), .C(stage0_r45_c38), .So(stage1_c83_s_fa0), .Co(stage1_c83_c_fa0));
    FA fa_802(.A(stage0_r46_c37), .B(stage0_r47_c36), .C(stage0_r48_c35), .So(stage1_c83_s_fa1), .Co(stage1_c83_c_fa1));
    FA fa_803(.A(stage0_r49_c34), .B(stage0_r50_c33), .C(stage0_r51_c32), .So(stage1_c83_s_fa2), .Co(stage1_c83_c_fa2));
    FA fa_804(.A(stage0_r52_c31), .B(stage0_r53_c30), .C(stage0_r54_c29), .So(stage1_c83_s_fa3), .Co(stage1_c83_c_fa3));
    FA fa_805(.A(stage0_r55_c28), .B(stage0_r56_c27), .C(stage0_r57_c26), .So(stage1_c83_s_fa4), .Co(stage1_c83_c_fa4));
    FA fa_806(.A(stage0_r58_c25), .B(stage0_r59_c24), .C(stage0_r60_c23), .So(stage1_c83_s_fa5), .Co(stage1_c83_c_fa5));
    FA fa_807(.A(stage0_r61_c22), .B(stage0_r62_c21), .C(stage0_r63_c20), .So(stage1_c83_s_fa6), .Co(stage1_c83_c_fa6));
    FA fa_808(.A(stage0_r64_c19), .B(stage0_r65_c18), .C(stage0_r66_c17), .So(stage1_c83_s_fa7), .Co(stage1_c83_c_fa7));
    FA fa_809(.A(stage0_r67_c16), .B(stage0_r68_c15), .C(stage0_r69_c14), .So(stage1_c83_s_fa8), .Co(stage1_c83_c_fa8));
    HA ha_48(.A(stage0_r70_c13), .B(stage0_r71_c12), .So(stage1_c83_s_ha0), .Co(stage1_c83_c_ha0));
    FA fa_810(.A(stage0_r44_c40), .B(stage0_r45_c39), .C(stage0_r46_c38), .So(stage1_c84_s_fa0), .Co(stage1_c84_c_fa0));
    FA fa_811(.A(stage0_r47_c37), .B(stage0_r48_c36), .C(stage0_r49_c35), .So(stage1_c84_s_fa1), .Co(stage1_c84_c_fa1));
    FA fa_812(.A(stage0_r50_c34), .B(stage0_r51_c33), .C(stage0_r52_c32), .So(stage1_c84_s_fa2), .Co(stage1_c84_c_fa2));
    FA fa_813(.A(stage0_r53_c31), .B(stage0_r54_c30), .C(stage0_r55_c29), .So(stage1_c84_s_fa3), .Co(stage1_c84_c_fa3));
    FA fa_814(.A(stage0_r56_c28), .B(stage0_r57_c27), .C(stage0_r58_c26), .So(stage1_c84_s_fa4), .Co(stage1_c84_c_fa4));
    FA fa_815(.A(stage0_r59_c25), .B(stage0_r60_c24), .C(stage0_r61_c23), .So(stage1_c84_s_fa5), .Co(stage1_c84_c_fa5));
    FA fa_816(.A(stage0_r62_c22), .B(stage0_r63_c21), .C(stage0_r64_c20), .So(stage1_c84_s_fa6), .Co(stage1_c84_c_fa6));
    FA fa_817(.A(stage0_r65_c19), .B(stage0_r66_c18), .C(stage0_r67_c17), .So(stage1_c84_s_fa7), .Co(stage1_c84_c_fa7));
    FA fa_818(.A(stage0_r68_c16), .B(stage0_r69_c15), .C(stage0_r70_c14), .So(stage1_c84_s_fa8), .Co(stage1_c84_c_fa8));
    FA fa_819(.A(stage0_r45_c40), .B(stage0_r46_c39), .C(stage0_r47_c38), .So(stage1_c85_s_fa0), .Co(stage1_c85_c_fa0));
    FA fa_820(.A(stage0_r48_c37), .B(stage0_r49_c36), .C(stage0_r50_c35), .So(stage1_c85_s_fa1), .Co(stage1_c85_c_fa1));
    FA fa_821(.A(stage0_r51_c34), .B(stage0_r52_c33), .C(stage0_r53_c32), .So(stage1_c85_s_fa2), .Co(stage1_c85_c_fa2));
    FA fa_822(.A(stage0_r54_c31), .B(stage0_r55_c30), .C(stage0_r56_c29), .So(stage1_c85_s_fa3), .Co(stage1_c85_c_fa3));
    FA fa_823(.A(stage0_r57_c28), .B(stage0_r58_c27), .C(stage0_r59_c26), .So(stage1_c85_s_fa4), .Co(stage1_c85_c_fa4));
    FA fa_824(.A(stage0_r60_c25), .B(stage0_r61_c24), .C(stage0_r62_c23), .So(stage1_c85_s_fa5), .Co(stage1_c85_c_fa5));
    FA fa_825(.A(stage0_r63_c22), .B(stage0_r64_c21), .C(stage0_r65_c20), .So(stage1_c85_s_fa6), .Co(stage1_c85_c_fa6));
    FA fa_826(.A(stage0_r66_c19), .B(stage0_r67_c18), .C(stage0_r68_c17), .So(stage1_c85_s_fa7), .Co(stage1_c85_c_fa7));
    FA fa_827(.A(stage0_r69_c16), .B(stage0_r70_c15), .C(stage0_r71_c14), .So(stage1_c85_s_fa8), .Co(stage1_c85_c_fa8));
    FA fa_828(.A(stage0_r46_c40), .B(stage0_r47_c39), .C(stage0_r48_c38), .So(stage1_c86_s_fa0), .Co(stage1_c86_c_fa0));
    FA fa_829(.A(stage0_r49_c37), .B(stage0_r50_c36), .C(stage0_r51_c35), .So(stage1_c86_s_fa1), .Co(stage1_c86_c_fa1));
    FA fa_830(.A(stage0_r52_c34), .B(stage0_r53_c33), .C(stage0_r54_c32), .So(stage1_c86_s_fa2), .Co(stage1_c86_c_fa2));
    FA fa_831(.A(stage0_r55_c31), .B(stage0_r56_c30), .C(stage0_r57_c29), .So(stage1_c86_s_fa3), .Co(stage1_c86_c_fa3));
    FA fa_832(.A(stage0_r58_c28), .B(stage0_r59_c27), .C(stage0_r60_c26), .So(stage1_c86_s_fa4), .Co(stage1_c86_c_fa4));
    FA fa_833(.A(stage0_r61_c25), .B(stage0_r62_c24), .C(stage0_r63_c23), .So(stage1_c86_s_fa5), .Co(stage1_c86_c_fa5));
    FA fa_834(.A(stage0_r64_c22), .B(stage0_r65_c21), .C(stage0_r66_c20), .So(stage1_c86_s_fa6), .Co(stage1_c86_c_fa6));
    FA fa_835(.A(stage0_r67_c19), .B(stage0_r68_c18), .C(stage0_r69_c17), .So(stage1_c86_s_fa7), .Co(stage1_c86_c_fa7));
    HA ha_49(.A(stage0_r70_c16), .B(stage0_r71_c15), .So(stage1_c86_s_ha0), .Co(stage1_c86_c_ha0));
    FA fa_836(.A(stage0_r47_c40), .B(stage0_r48_c39), .C(stage0_r49_c38), .So(stage1_c87_s_fa0), .Co(stage1_c87_c_fa0));
    FA fa_837(.A(stage0_r50_c37), .B(stage0_r51_c36), .C(stage0_r52_c35), .So(stage1_c87_s_fa1), .Co(stage1_c87_c_fa1));
    FA fa_838(.A(stage0_r53_c34), .B(stage0_r54_c33), .C(stage0_r55_c32), .So(stage1_c87_s_fa2), .Co(stage1_c87_c_fa2));
    FA fa_839(.A(stage0_r56_c31), .B(stage0_r57_c30), .C(stage0_r58_c29), .So(stage1_c87_s_fa3), .Co(stage1_c87_c_fa3));
    FA fa_840(.A(stage0_r59_c28), .B(stage0_r60_c27), .C(stage0_r61_c26), .So(stage1_c87_s_fa4), .Co(stage1_c87_c_fa4));
    FA fa_841(.A(stage0_r62_c25), .B(stage0_r63_c24), .C(stage0_r64_c23), .So(stage1_c87_s_fa5), .Co(stage1_c87_c_fa5));
    FA fa_842(.A(stage0_r65_c22), .B(stage0_r66_c21), .C(stage0_r67_c20), .So(stage1_c87_s_fa6), .Co(stage1_c87_c_fa6));
    FA fa_843(.A(stage0_r68_c19), .B(stage0_r69_c18), .C(stage0_r70_c17), .So(stage1_c87_s_fa7), .Co(stage1_c87_c_fa7));
    FA fa_844(.A(stage0_r48_c40), .B(stage0_r49_c39), .C(stage0_r50_c38), .So(stage1_c88_s_fa0), .Co(stage1_c88_c_fa0));
    FA fa_845(.A(stage0_r51_c37), .B(stage0_r52_c36), .C(stage0_r53_c35), .So(stage1_c88_s_fa1), .Co(stage1_c88_c_fa1));
    FA fa_846(.A(stage0_r54_c34), .B(stage0_r55_c33), .C(stage0_r56_c32), .So(stage1_c88_s_fa2), .Co(stage1_c88_c_fa2));
    FA fa_847(.A(stage0_r57_c31), .B(stage0_r58_c30), .C(stage0_r59_c29), .So(stage1_c88_s_fa3), .Co(stage1_c88_c_fa3));
    FA fa_848(.A(stage0_r60_c28), .B(stage0_r61_c27), .C(stage0_r62_c26), .So(stage1_c88_s_fa4), .Co(stage1_c88_c_fa4));
    FA fa_849(.A(stage0_r63_c25), .B(stage0_r64_c24), .C(stage0_r65_c23), .So(stage1_c88_s_fa5), .Co(stage1_c88_c_fa5));
    FA fa_850(.A(stage0_r66_c22), .B(stage0_r67_c21), .C(stage0_r68_c20), .So(stage1_c88_s_fa6), .Co(stage1_c88_c_fa6));
    FA fa_851(.A(stage0_r69_c19), .B(stage0_r70_c18), .C(stage0_r71_c17), .So(stage1_c88_s_fa7), .Co(stage1_c88_c_fa7));
    FA fa_852(.A(stage0_r49_c40), .B(stage0_r50_c39), .C(stage0_r51_c38), .So(stage1_c89_s_fa0), .Co(stage1_c89_c_fa0));
    FA fa_853(.A(stage0_r52_c37), .B(stage0_r53_c36), .C(stage0_r54_c35), .So(stage1_c89_s_fa1), .Co(stage1_c89_c_fa1));
    FA fa_854(.A(stage0_r55_c34), .B(stage0_r56_c33), .C(stage0_r57_c32), .So(stage1_c89_s_fa2), .Co(stage1_c89_c_fa2));
    FA fa_855(.A(stage0_r58_c31), .B(stage0_r59_c30), .C(stage0_r60_c29), .So(stage1_c89_s_fa3), .Co(stage1_c89_c_fa3));
    FA fa_856(.A(stage0_r61_c28), .B(stage0_r62_c27), .C(stage0_r63_c26), .So(stage1_c89_s_fa4), .Co(stage1_c89_c_fa4));
    FA fa_857(.A(stage0_r64_c25), .B(stage0_r65_c24), .C(stage0_r66_c23), .So(stage1_c89_s_fa5), .Co(stage1_c89_c_fa5));
    FA fa_858(.A(stage0_r67_c22), .B(stage0_r68_c21), .C(stage0_r69_c20), .So(stage1_c89_s_fa6), .Co(stage1_c89_c_fa6));
    HA ha_50(.A(stage0_r70_c19), .B(stage0_r71_c18), .So(stage1_c89_s_ha0), .Co(stage1_c89_c_ha0));
    FA fa_859(.A(stage0_r50_c40), .B(stage0_r51_c39), .C(stage0_r52_c38), .So(stage1_c90_s_fa0), .Co(stage1_c90_c_fa0));
    FA fa_860(.A(stage0_r53_c37), .B(stage0_r54_c36), .C(stage0_r55_c35), .So(stage1_c90_s_fa1), .Co(stage1_c90_c_fa1));
    FA fa_861(.A(stage0_r56_c34), .B(stage0_r57_c33), .C(stage0_r58_c32), .So(stage1_c90_s_fa2), .Co(stage1_c90_c_fa2));
    FA fa_862(.A(stage0_r59_c31), .B(stage0_r60_c30), .C(stage0_r61_c29), .So(stage1_c90_s_fa3), .Co(stage1_c90_c_fa3));
    FA fa_863(.A(stage0_r62_c28), .B(stage0_r63_c27), .C(stage0_r64_c26), .So(stage1_c90_s_fa4), .Co(stage1_c90_c_fa4));
    FA fa_864(.A(stage0_r65_c25), .B(stage0_r66_c24), .C(stage0_r67_c23), .So(stage1_c90_s_fa5), .Co(stage1_c90_c_fa5));
    FA fa_865(.A(stage0_r68_c22), .B(stage0_r69_c21), .C(stage0_r70_c20), .So(stage1_c90_s_fa6), .Co(stage1_c90_c_fa6));
    FA fa_866(.A(stage0_r51_c40), .B(stage0_r52_c39), .C(stage0_r53_c38), .So(stage1_c91_s_fa0), .Co(stage1_c91_c_fa0));
    FA fa_867(.A(stage0_r54_c37), .B(stage0_r55_c36), .C(stage0_r56_c35), .So(stage1_c91_s_fa1), .Co(stage1_c91_c_fa1));
    FA fa_868(.A(stage0_r57_c34), .B(stage0_r58_c33), .C(stage0_r59_c32), .So(stage1_c91_s_fa2), .Co(stage1_c91_c_fa2));
    FA fa_869(.A(stage0_r60_c31), .B(stage0_r61_c30), .C(stage0_r62_c29), .So(stage1_c91_s_fa3), .Co(stage1_c91_c_fa3));
    FA fa_870(.A(stage0_r63_c28), .B(stage0_r64_c27), .C(stage0_r65_c26), .So(stage1_c91_s_fa4), .Co(stage1_c91_c_fa4));
    FA fa_871(.A(stage0_r66_c25), .B(stage0_r67_c24), .C(stage0_r68_c23), .So(stage1_c91_s_fa5), .Co(stage1_c91_c_fa5));
    FA fa_872(.A(stage0_r69_c22), .B(stage0_r70_c21), .C(stage0_r71_c20), .So(stage1_c91_s_fa6), .Co(stage1_c91_c_fa6));
    FA fa_873(.A(stage0_r52_c40), .B(stage0_r53_c39), .C(stage0_r54_c38), .So(stage1_c92_s_fa0), .Co(stage1_c92_c_fa0));
    FA fa_874(.A(stage0_r55_c37), .B(stage0_r56_c36), .C(stage0_r57_c35), .So(stage1_c92_s_fa1), .Co(stage1_c92_c_fa1));
    FA fa_875(.A(stage0_r58_c34), .B(stage0_r59_c33), .C(stage0_r60_c32), .So(stage1_c92_s_fa2), .Co(stage1_c92_c_fa2));
    FA fa_876(.A(stage0_r61_c31), .B(stage0_r62_c30), .C(stage0_r63_c29), .So(stage1_c92_s_fa3), .Co(stage1_c92_c_fa3));
    FA fa_877(.A(stage0_r64_c28), .B(stage0_r65_c27), .C(stage0_r66_c26), .So(stage1_c92_s_fa4), .Co(stage1_c92_c_fa4));
    FA fa_878(.A(stage0_r67_c25), .B(stage0_r68_c24), .C(stage0_r69_c23), .So(stage1_c92_s_fa5), .Co(stage1_c92_c_fa5));
    HA ha_51(.A(stage0_r70_c22), .B(stage0_r71_c21), .So(stage1_c92_s_ha0), .Co(stage1_c92_c_ha0));
    FA fa_879(.A(stage0_r53_c40), .B(stage0_r54_c39), .C(stage0_r55_c38), .So(stage1_c93_s_fa0), .Co(stage1_c93_c_fa0));
    FA fa_880(.A(stage0_r56_c37), .B(stage0_r57_c36), .C(stage0_r58_c35), .So(stage1_c93_s_fa1), .Co(stage1_c93_c_fa1));
    FA fa_881(.A(stage0_r59_c34), .B(stage0_r60_c33), .C(stage0_r61_c32), .So(stage1_c93_s_fa2), .Co(stage1_c93_c_fa2));
    FA fa_882(.A(stage0_r62_c31), .B(stage0_r63_c30), .C(stage0_r64_c29), .So(stage1_c93_s_fa3), .Co(stage1_c93_c_fa3));
    FA fa_883(.A(stage0_r65_c28), .B(stage0_r66_c27), .C(stage0_r67_c26), .So(stage1_c93_s_fa4), .Co(stage1_c93_c_fa4));
    FA fa_884(.A(stage0_r68_c25), .B(stage0_r69_c24), .C(stage0_r70_c23), .So(stage1_c93_s_fa5), .Co(stage1_c93_c_fa5));
    FA fa_885(.A(stage0_r54_c40), .B(stage0_r55_c39), .C(stage0_r56_c38), .So(stage1_c94_s_fa0), .Co(stage1_c94_c_fa0));
    FA fa_886(.A(stage0_r57_c37), .B(stage0_r58_c36), .C(stage0_r59_c35), .So(stage1_c94_s_fa1), .Co(stage1_c94_c_fa1));
    FA fa_887(.A(stage0_r60_c34), .B(stage0_r61_c33), .C(stage0_r62_c32), .So(stage1_c94_s_fa2), .Co(stage1_c94_c_fa2));
    FA fa_888(.A(stage0_r63_c31), .B(stage0_r64_c30), .C(stage0_r65_c29), .So(stage1_c94_s_fa3), .Co(stage1_c94_c_fa3));
    FA fa_889(.A(stage0_r66_c28), .B(stage0_r67_c27), .C(stage0_r68_c26), .So(stage1_c94_s_fa4), .Co(stage1_c94_c_fa4));
    FA fa_890(.A(stage0_r69_c25), .B(stage0_r70_c24), .C(stage0_r71_c23), .So(stage1_c94_s_fa5), .Co(stage1_c94_c_fa5));
    FA fa_891(.A(stage0_r55_c40), .B(stage0_r56_c39), .C(stage0_r57_c38), .So(stage1_c95_s_fa0), .Co(stage1_c95_c_fa0));
    FA fa_892(.A(stage0_r58_c37), .B(stage0_r59_c36), .C(stage0_r60_c35), .So(stage1_c95_s_fa1), .Co(stage1_c95_c_fa1));
    FA fa_893(.A(stage0_r61_c34), .B(stage0_r62_c33), .C(stage0_r63_c32), .So(stage1_c95_s_fa2), .Co(stage1_c95_c_fa2));
    FA fa_894(.A(stage0_r64_c31), .B(stage0_r65_c30), .C(stage0_r66_c29), .So(stage1_c95_s_fa3), .Co(stage1_c95_c_fa3));
    FA fa_895(.A(stage0_r67_c28), .B(stage0_r68_c27), .C(stage0_r69_c26), .So(stage1_c95_s_fa4), .Co(stage1_c95_c_fa4));
    HA ha_52(.A(stage0_r70_c25), .B(stage0_r71_c24), .So(stage1_c95_s_ha0), .Co(stage1_c95_c_ha0));
    FA fa_896(.A(stage0_r56_c40), .B(stage0_r57_c39), .C(stage0_r58_c38), .So(stage1_c96_s_fa0), .Co(stage1_c96_c_fa0));
    FA fa_897(.A(stage0_r59_c37), .B(stage0_r60_c36), .C(stage0_r61_c35), .So(stage1_c96_s_fa1), .Co(stage1_c96_c_fa1));
    FA fa_898(.A(stage0_r62_c34), .B(stage0_r63_c33), .C(stage0_r64_c32), .So(stage1_c96_s_fa2), .Co(stage1_c96_c_fa2));
    FA fa_899(.A(stage0_r65_c31), .B(stage0_r66_c30), .C(stage0_r67_c29), .So(stage1_c96_s_fa3), .Co(stage1_c96_c_fa3));
    FA fa_900(.A(stage0_r68_c28), .B(stage0_r69_c27), .C(stage0_r70_c26), .So(stage1_c96_s_fa4), .Co(stage1_c96_c_fa4));
    FA fa_901(.A(stage0_r57_c40), .B(stage0_r58_c39), .C(stage0_r59_c38), .So(stage1_c97_s_fa0), .Co(stage1_c97_c_fa0));
    FA fa_902(.A(stage0_r60_c37), .B(stage0_r61_c36), .C(stage0_r62_c35), .So(stage1_c97_s_fa1), .Co(stage1_c97_c_fa1));
    FA fa_903(.A(stage0_r63_c34), .B(stage0_r64_c33), .C(stage0_r65_c32), .So(stage1_c97_s_fa2), .Co(stage1_c97_c_fa2));
    FA fa_904(.A(stage0_r66_c31), .B(stage0_r67_c30), .C(stage0_r68_c29), .So(stage1_c97_s_fa3), .Co(stage1_c97_c_fa3));
    FA fa_905(.A(stage0_r69_c28), .B(stage0_r70_c27), .C(stage0_r71_c26), .So(stage1_c97_s_fa4), .Co(stage1_c97_c_fa4));
    FA fa_906(.A(stage0_r58_c40), .B(stage0_r59_c39), .C(stage0_r60_c38), .So(stage1_c98_s_fa0), .Co(stage1_c98_c_fa0));
    FA fa_907(.A(stage0_r61_c37), .B(stage0_r62_c36), .C(stage0_r63_c35), .So(stage1_c98_s_fa1), .Co(stage1_c98_c_fa1));
    FA fa_908(.A(stage0_r64_c34), .B(stage0_r65_c33), .C(stage0_r66_c32), .So(stage1_c98_s_fa2), .Co(stage1_c98_c_fa2));
    FA fa_909(.A(stage0_r67_c31), .B(stage0_r68_c30), .C(stage0_r69_c29), .So(stage1_c98_s_fa3), .Co(stage1_c98_c_fa3));
    HA ha_53(.A(stage0_r70_c28), .B(stage0_r71_c27), .So(stage1_c98_s_ha0), .Co(stage1_c98_c_ha0));
    FA fa_910(.A(stage0_r59_c40), .B(stage0_r60_c39), .C(stage0_r61_c38), .So(stage1_c99_s_fa0), .Co(stage1_c99_c_fa0));
    FA fa_911(.A(stage0_r62_c37), .B(stage0_r63_c36), .C(stage0_r64_c35), .So(stage1_c99_s_fa1), .Co(stage1_c99_c_fa1));
    FA fa_912(.A(stage0_r65_c34), .B(stage0_r66_c33), .C(stage0_r67_c32), .So(stage1_c99_s_fa2), .Co(stage1_c99_c_fa2));
    FA fa_913(.A(stage0_r68_c31), .B(stage0_r69_c30), .C(stage0_r70_c29), .So(stage1_c99_s_fa3), .Co(stage1_c99_c_fa3));
    FA fa_914(.A(stage0_r60_c40), .B(stage0_r61_c39), .C(stage0_r62_c38), .So(stage1_c100_s_fa0), .Co(stage1_c100_c_fa0));
    FA fa_915(.A(stage0_r63_c37), .B(stage0_r64_c36), .C(stage0_r65_c35), .So(stage1_c100_s_fa1), .Co(stage1_c100_c_fa1));
    FA fa_916(.A(stage0_r66_c34), .B(stage0_r67_c33), .C(stage0_r68_c32), .So(stage1_c100_s_fa2), .Co(stage1_c100_c_fa2));
    FA fa_917(.A(stage0_r69_c31), .B(stage0_r70_c30), .C(stage0_r71_c29), .So(stage1_c100_s_fa3), .Co(stage1_c100_c_fa3));
    FA fa_918(.A(stage0_r61_c40), .B(stage0_r62_c39), .C(stage0_r63_c38), .So(stage1_c101_s_fa0), .Co(stage1_c101_c_fa0));
    FA fa_919(.A(stage0_r64_c37), .B(stage0_r65_c36), .C(stage0_r66_c35), .So(stage1_c101_s_fa1), .Co(stage1_c101_c_fa1));
    FA fa_920(.A(stage0_r67_c34), .B(stage0_r68_c33), .C(stage0_r69_c32), .So(stage1_c101_s_fa2), .Co(stage1_c101_c_fa2));
    HA ha_54(.A(stage0_r70_c31), .B(stage0_r71_c30), .So(stage1_c101_s_ha0), .Co(stage1_c101_c_ha0));
    FA fa_921(.A(stage0_r62_c40), .B(stage0_r63_c39), .C(stage0_r64_c38), .So(stage1_c102_s_fa0), .Co(stage1_c102_c_fa0));
    FA fa_922(.A(stage0_r65_c37), .B(stage0_r66_c36), .C(stage0_r67_c35), .So(stage1_c102_s_fa1), .Co(stage1_c102_c_fa1));
    FA fa_923(.A(stage0_r68_c34), .B(stage0_r69_c33), .C(stage0_r70_c32), .So(stage1_c102_s_fa2), .Co(stage1_c102_c_fa2));
    FA fa_924(.A(stage0_r63_c40), .B(stage0_r64_c39), .C(stage0_r65_c38), .So(stage1_c103_s_fa0), .Co(stage1_c103_c_fa0));
    FA fa_925(.A(stage0_r66_c37), .B(stage0_r67_c36), .C(stage0_r68_c35), .So(stage1_c103_s_fa1), .Co(stage1_c103_c_fa1));
    FA fa_926(.A(stage0_r69_c34), .B(stage0_r70_c33), .C(stage0_r71_c32), .So(stage1_c103_s_fa2), .Co(stage1_c103_c_fa2));
    FA fa_927(.A(stage0_r64_c40), .B(stage0_r65_c39), .C(stage0_r66_c38), .So(stage1_c104_s_fa0), .Co(stage1_c104_c_fa0));
    FA fa_928(.A(stage0_r67_c37), .B(stage0_r68_c36), .C(stage0_r69_c35), .So(stage1_c104_s_fa1), .Co(stage1_c104_c_fa1));
    HA ha_55(.A(stage0_r70_c34), .B(stage0_r71_c33), .So(stage1_c104_s_ha0), .Co(stage1_c104_c_ha0));
    FA fa_929(.A(stage0_r65_c40), .B(stage0_r66_c39), .C(stage0_r67_c38), .So(stage1_c105_s_fa0), .Co(stage1_c105_c_fa0));
    FA fa_930(.A(stage0_r68_c37), .B(stage0_r69_c36), .C(stage0_r70_c35), .So(stage1_c105_s_fa1), .Co(stage1_c105_c_fa1));
    FA fa_931(.A(stage0_r66_c40), .B(stage0_r67_c39), .C(stage0_r68_c38), .So(stage1_c106_s_fa0), .Co(stage1_c106_c_fa0));
    FA fa_932(.A(stage0_r69_c37), .B(stage0_r70_c36), .C(stage0_r71_c35), .So(stage1_c106_s_fa1), .Co(stage1_c106_c_fa1));
    FA fa_933(.A(stage0_r67_c40), .B(stage0_r68_c39), .C(stage0_r69_c38), .So(stage1_c107_s_fa0), .Co(stage1_c107_c_fa0));
    HA ha_56(.A(stage0_r70_c37), .B(stage0_r71_c36), .So(stage1_c107_s_ha0), .Co(stage1_c107_c_ha0));
    FA fa_934(.A(stage0_r68_c40), .B(stage0_r69_c39), .C(stage0_r70_c38), .So(stage1_c108_s_fa0), .Co(stage1_c108_c_fa0));
    FA fa_935(.A(stage0_r69_c40), .B(stage0_r70_c39), .C(stage0_r71_c38), .So(stage1_c109_s_fa0), .Co(stage1_c109_c_fa0));
    HA ha_57(.A(stage0_r70_c40), .B(stage0_r71_c39), .So(stage1_c110_s_ha0), .Co(stage1_c110_c_ha0));
    HA ha_58(.A(stage1_c1_c_ha0), .B(stage1_c2_s_fa0), .So(stage2_c2_s_ha0), .Co(stage2_c2_c_ha0));
    FA fa_936(.A(stage1_c2_c_fa0), .B(stage1_c3_s_fa0), .C(stage0_r3_c0), .So(stage2_c3_s_fa0), .Co(stage2_c3_c_fa0));
    FA fa_937(.A(stage1_c3_c_fa0), .B(stage1_c4_s_fa0), .C(stage1_c4_s_ha0), .So(stage2_c4_s_fa0), .Co(stage2_c4_c_fa0));
    FA fa_938(.A(stage1_c4_c_fa0), .B(stage1_c4_c_ha0), .C(stage1_c5_s_fa0), .So(stage2_c5_s_fa0), .Co(stage2_c5_c_fa0));
    FA fa_939(.A(stage1_c5_c_fa0), .B(stage1_c5_c_fa1), .C(stage1_c6_s_fa0), .So(stage2_c6_s_fa0), .Co(stage2_c6_c_fa0));
    HA ha_59(.A(stage1_c6_s_fa1), .B(stage0_r6_c0), .So(stage2_c6_s_ha0), .Co(stage2_c6_c_ha0));
    FA fa_940(.A(stage1_c6_c_fa0), .B(stage1_c6_c_fa1), .C(stage1_c7_s_fa0), .So(stage2_c7_s_fa0), .Co(stage2_c7_c_fa0));
    HA ha_60(.A(stage1_c7_s_fa1), .B(stage1_c7_s_ha0), .So(stage2_c7_s_ha0), .Co(stage2_c7_c_ha0));
    FA fa_941(.A(stage1_c7_c_fa0), .B(stage1_c7_c_fa1), .C(stage1_c7_c_ha0), .So(stage2_c8_s_fa0), .Co(stage2_c8_c_fa0));
    FA fa_942(.A(stage1_c8_s_fa0), .B(stage1_c8_s_fa1), .C(stage1_c8_s_fa2), .So(stage2_c8_s_fa1), .Co(stage2_c8_c_fa1));
    FA fa_943(.A(stage1_c8_c_fa0), .B(stage1_c8_c_fa1), .C(stage1_c8_c_fa2), .So(stage2_c9_s_fa0), .Co(stage2_c9_c_fa0));
    FA fa_944(.A(stage1_c9_s_fa0), .B(stage1_c9_s_fa1), .C(stage1_c9_s_fa2), .So(stage2_c9_s_fa1), .Co(stage2_c9_c_fa1));
    FA fa_945(.A(stage1_c9_c_fa0), .B(stage1_c9_c_fa1), .C(stage1_c9_c_fa2), .So(stage2_c10_s_fa0), .Co(stage2_c10_c_fa0));
    FA fa_946(.A(stage1_c10_s_fa0), .B(stage1_c10_s_fa1), .C(stage1_c10_s_fa2), .So(stage2_c10_s_fa1), .Co(stage2_c10_c_fa1));
    FA fa_947(.A(stage1_c10_c_fa0), .B(stage1_c10_c_fa1), .C(stage1_c10_c_fa2), .So(stage2_c11_s_fa0), .Co(stage2_c11_c_fa0));
    FA fa_948(.A(stage1_c10_c_ha0), .B(stage1_c11_s_fa0), .C(stage1_c11_s_fa1), .So(stage2_c11_s_fa1), .Co(stage2_c11_c_fa1));
    HA ha_61(.A(stage1_c11_s_fa2), .B(stage1_c11_s_fa3), .So(stage2_c11_s_ha0), .Co(stage2_c11_c_ha0));
    FA fa_949(.A(stage1_c11_c_fa0), .B(stage1_c11_c_fa1), .C(stage1_c11_c_fa2), .So(stage2_c12_s_fa0), .Co(stage2_c12_c_fa0));
    FA fa_950(.A(stage1_c11_c_fa3), .B(stage1_c12_s_fa0), .C(stage1_c12_s_fa1), .So(stage2_c12_s_fa1), .Co(stage2_c12_c_fa1));
    FA fa_951(.A(stage1_c12_s_fa2), .B(stage1_c12_s_fa3), .C(stage0_r12_c0), .So(stage2_c12_s_fa2), .Co(stage2_c12_c_fa2));
    FA fa_952(.A(stage1_c12_c_fa0), .B(stage1_c12_c_fa1), .C(stage1_c12_c_fa2), .So(stage2_c13_s_fa0), .Co(stage2_c13_c_fa0));
    FA fa_953(.A(stage1_c12_c_fa3), .B(stage1_c13_s_fa0), .C(stage1_c13_s_fa1), .So(stage2_c13_s_fa1), .Co(stage2_c13_c_fa1));
    FA fa_954(.A(stage1_c13_s_fa2), .B(stage1_c13_s_fa3), .C(stage1_c13_s_ha0), .So(stage2_c13_s_fa2), .Co(stage2_c13_c_fa2));
    FA fa_955(.A(stage1_c13_c_fa0), .B(stage1_c13_c_fa1), .C(stage1_c13_c_fa2), .So(stage2_c14_s_fa0), .Co(stage2_c14_c_fa0));
    FA fa_956(.A(stage1_c13_c_fa3), .B(stage1_c13_c_ha0), .C(stage1_c14_s_fa0), .So(stage2_c14_s_fa1), .Co(stage2_c14_c_fa1));
    FA fa_957(.A(stage1_c14_s_fa1), .B(stage1_c14_s_fa2), .C(stage1_c14_s_fa3), .So(stage2_c14_s_fa2), .Co(stage2_c14_c_fa2));
    FA fa_958(.A(stage1_c14_c_fa0), .B(stage1_c14_c_fa1), .C(stage1_c14_c_fa2), .So(stage2_c15_s_fa0), .Co(stage2_c15_c_fa0));
    FA fa_959(.A(stage1_c14_c_fa3), .B(stage1_c14_c_fa4), .C(stage1_c15_s_fa0), .So(stage2_c15_s_fa1), .Co(stage2_c15_c_fa1));
    FA fa_960(.A(stage1_c15_s_fa1), .B(stage1_c15_s_fa2), .C(stage1_c15_s_fa3), .So(stage2_c15_s_fa2), .Co(stage2_c15_c_fa2));
    HA ha_62(.A(stage1_c15_s_fa4), .B(stage0_r15_c0), .So(stage2_c15_s_ha0), .Co(stage2_c15_c_ha0));
    FA fa_961(.A(stage1_c15_c_fa0), .B(stage1_c15_c_fa1), .C(stage1_c15_c_fa2), .So(stage2_c16_s_fa0), .Co(stage2_c16_c_fa0));
    FA fa_962(.A(stage1_c15_c_fa3), .B(stage1_c15_c_fa4), .C(stage1_c16_s_fa0), .So(stage2_c16_s_fa1), .Co(stage2_c16_c_fa1));
    FA fa_963(.A(stage1_c16_s_fa1), .B(stage1_c16_s_fa2), .C(stage1_c16_s_fa3), .So(stage2_c16_s_fa2), .Co(stage2_c16_c_fa2));
    HA ha_63(.A(stage1_c16_s_fa4), .B(stage1_c16_s_ha0), .So(stage2_c16_s_ha0), .Co(stage2_c16_c_ha0));
    FA fa_964(.A(stage1_c16_c_fa0), .B(stage1_c16_c_fa1), .C(stage1_c16_c_fa2), .So(stage2_c17_s_fa0), .Co(stage2_c17_c_fa0));
    FA fa_965(.A(stage1_c16_c_fa3), .B(stage1_c16_c_fa4), .C(stage1_c16_c_ha0), .So(stage2_c17_s_fa1), .Co(stage2_c17_c_fa1));
    FA fa_966(.A(stage1_c17_s_fa0), .B(stage1_c17_s_fa1), .C(stage1_c17_s_fa2), .So(stage2_c17_s_fa2), .Co(stage2_c17_c_fa2));
    FA fa_967(.A(stage1_c17_s_fa3), .B(stage1_c17_s_fa4), .C(stage1_c17_s_fa5), .So(stage2_c17_s_fa3), .Co(stage2_c17_c_fa3));
    FA fa_968(.A(stage1_c17_c_fa0), .B(stage1_c17_c_fa1), .C(stage1_c17_c_fa2), .So(stage2_c18_s_fa0), .Co(stage2_c18_c_fa0));
    FA fa_969(.A(stage1_c17_c_fa3), .B(stage1_c17_c_fa4), .C(stage1_c17_c_fa5), .So(stage2_c18_s_fa1), .Co(stage2_c18_c_fa1));
    FA fa_970(.A(stage1_c18_s_fa0), .B(stage1_c18_s_fa1), .C(stage1_c18_s_fa2), .So(stage2_c18_s_fa2), .Co(stage2_c18_c_fa2));
    FA fa_971(.A(stage1_c18_s_fa3), .B(stage1_c18_s_fa4), .C(stage1_c18_s_fa5), .So(stage2_c18_s_fa3), .Co(stage2_c18_c_fa3));
    FA fa_972(.A(stage1_c18_c_fa0), .B(stage1_c18_c_fa1), .C(stage1_c18_c_fa2), .So(stage2_c19_s_fa0), .Co(stage2_c19_c_fa0));
    FA fa_973(.A(stage1_c18_c_fa3), .B(stage1_c18_c_fa4), .C(stage1_c18_c_fa5), .So(stage2_c19_s_fa1), .Co(stage2_c19_c_fa1));
    FA fa_974(.A(stage1_c19_s_fa0), .B(stage1_c19_s_fa1), .C(stage1_c19_s_fa2), .So(stage2_c19_s_fa2), .Co(stage2_c19_c_fa2));
    FA fa_975(.A(stage1_c19_s_fa3), .B(stage1_c19_s_fa4), .C(stage1_c19_s_fa5), .So(stage2_c19_s_fa3), .Co(stage2_c19_c_fa3));
    FA fa_976(.A(stage1_c19_c_fa0), .B(stage1_c19_c_fa1), .C(stage1_c19_c_fa2), .So(stage2_c20_s_fa0), .Co(stage2_c20_c_fa0));
    FA fa_977(.A(stage1_c19_c_fa3), .B(stage1_c19_c_fa4), .C(stage1_c19_c_fa5), .So(stage2_c20_s_fa1), .Co(stage2_c20_c_fa1));
    FA fa_978(.A(stage1_c19_c_ha0), .B(stage1_c20_s_fa0), .C(stage1_c20_s_fa1), .So(stage2_c20_s_fa2), .Co(stage2_c20_c_fa2));
    FA fa_979(.A(stage1_c20_s_fa2), .B(stage1_c20_s_fa3), .C(stage1_c20_s_fa4), .So(stage2_c20_s_fa3), .Co(stage2_c20_c_fa3));
    HA ha_64(.A(stage1_c20_s_fa5), .B(stage1_c20_s_fa6), .So(stage2_c20_s_ha0), .Co(stage2_c20_c_ha0));
    FA fa_980(.A(stage1_c20_c_fa0), .B(stage1_c20_c_fa1), .C(stage1_c20_c_fa2), .So(stage2_c21_s_fa0), .Co(stage2_c21_c_fa0));
    FA fa_981(.A(stage1_c20_c_fa3), .B(stage1_c20_c_fa4), .C(stage1_c20_c_fa5), .So(stage2_c21_s_fa1), .Co(stage2_c21_c_fa1));
    FA fa_982(.A(stage1_c20_c_fa6), .B(stage1_c21_s_fa0), .C(stage1_c21_s_fa1), .So(stage2_c21_s_fa2), .Co(stage2_c21_c_fa2));
    FA fa_983(.A(stage1_c21_s_fa2), .B(stage1_c21_s_fa3), .C(stage1_c21_s_fa4), .So(stage2_c21_s_fa3), .Co(stage2_c21_c_fa3));
    FA fa_984(.A(stage1_c21_s_fa5), .B(stage1_c21_s_fa6), .C(stage0_r21_c0), .So(stage2_c21_s_fa4), .Co(stage2_c21_c_fa4));
    FA fa_985(.A(stage1_c21_c_fa0), .B(stage1_c21_c_fa1), .C(stage1_c21_c_fa2), .So(stage2_c22_s_fa0), .Co(stage2_c22_c_fa0));
    FA fa_986(.A(stage1_c21_c_fa3), .B(stage1_c21_c_fa4), .C(stage1_c21_c_fa5), .So(stage2_c22_s_fa1), .Co(stage2_c22_c_fa1));
    FA fa_987(.A(stage1_c21_c_fa6), .B(stage1_c22_s_fa0), .C(stage1_c22_s_fa1), .So(stage2_c22_s_fa2), .Co(stage2_c22_c_fa2));
    FA fa_988(.A(stage1_c22_s_fa2), .B(stage1_c22_s_fa3), .C(stage1_c22_s_fa4), .So(stage2_c22_s_fa3), .Co(stage2_c22_c_fa3));
    FA fa_989(.A(stage1_c22_s_fa5), .B(stage1_c22_s_fa6), .C(stage1_c22_s_ha0), .So(stage2_c22_s_fa4), .Co(stage2_c22_c_fa4));
    FA fa_990(.A(stage1_c22_c_fa0), .B(stage1_c22_c_fa1), .C(stage1_c22_c_fa2), .So(stage2_c23_s_fa0), .Co(stage2_c23_c_fa0));
    FA fa_991(.A(stage1_c22_c_fa3), .B(stage1_c22_c_fa4), .C(stage1_c22_c_fa5), .So(stage2_c23_s_fa1), .Co(stage2_c23_c_fa1));
    FA fa_992(.A(stage1_c22_c_fa6), .B(stage1_c22_c_ha0), .C(stage1_c23_s_fa0), .So(stage2_c23_s_fa2), .Co(stage2_c23_c_fa2));
    FA fa_993(.A(stage1_c23_s_fa1), .B(stage1_c23_s_fa2), .C(stage1_c23_s_fa3), .So(stage2_c23_s_fa3), .Co(stage2_c23_c_fa3));
    FA fa_994(.A(stage1_c23_s_fa4), .B(stage1_c23_s_fa5), .C(stage1_c23_s_fa6), .So(stage2_c23_s_fa4), .Co(stage2_c23_c_fa4));
    FA fa_995(.A(stage1_c23_c_fa0), .B(stage1_c23_c_fa1), .C(stage1_c23_c_fa2), .So(stage2_c24_s_fa0), .Co(stage2_c24_c_fa0));
    FA fa_996(.A(stage1_c23_c_fa3), .B(stage1_c23_c_fa4), .C(stage1_c23_c_fa5), .So(stage2_c24_s_fa1), .Co(stage2_c24_c_fa1));
    FA fa_997(.A(stage1_c23_c_fa6), .B(stage1_c23_c_fa7), .C(stage1_c24_s_fa0), .So(stage2_c24_s_fa2), .Co(stage2_c24_c_fa2));
    FA fa_998(.A(stage1_c24_s_fa1), .B(stage1_c24_s_fa2), .C(stage1_c24_s_fa3), .So(stage2_c24_s_fa3), .Co(stage2_c24_c_fa3));
    FA fa_999(.A(stage1_c24_s_fa4), .B(stage1_c24_s_fa5), .C(stage1_c24_s_fa6), .So(stage2_c24_s_fa4), .Co(stage2_c24_c_fa4));
    HA ha_65(.A(stage1_c24_s_fa7), .B(stage0_r24_c0), .So(stage2_c24_s_ha0), .Co(stage2_c24_c_ha0));
    FA fa_1000(.A(stage1_c24_c_fa0), .B(stage1_c24_c_fa1), .C(stage1_c24_c_fa2), .So(stage2_c25_s_fa0), .Co(stage2_c25_c_fa0));
    FA fa_1001(.A(stage1_c24_c_fa3), .B(stage1_c24_c_fa4), .C(stage1_c24_c_fa5), .So(stage2_c25_s_fa1), .Co(stage2_c25_c_fa1));
    FA fa_1002(.A(stage1_c24_c_fa6), .B(stage1_c24_c_fa7), .C(stage1_c25_s_fa0), .So(stage2_c25_s_fa2), .Co(stage2_c25_c_fa2));
    FA fa_1003(.A(stage1_c25_s_fa1), .B(stage1_c25_s_fa2), .C(stage1_c25_s_fa3), .So(stage2_c25_s_fa3), .Co(stage2_c25_c_fa3));
    FA fa_1004(.A(stage1_c25_s_fa4), .B(stage1_c25_s_fa5), .C(stage1_c25_s_fa6), .So(stage2_c25_s_fa4), .Co(stage2_c25_c_fa4));
    HA ha_66(.A(stage1_c25_s_fa7), .B(stage1_c25_s_ha0), .So(stage2_c25_s_ha0), .Co(stage2_c25_c_ha0));
    FA fa_1005(.A(stage1_c25_c_fa0), .B(stage1_c25_c_fa1), .C(stage1_c25_c_fa2), .So(stage2_c26_s_fa0), .Co(stage2_c26_c_fa0));
    FA fa_1006(.A(stage1_c25_c_fa3), .B(stage1_c25_c_fa4), .C(stage1_c25_c_fa5), .So(stage2_c26_s_fa1), .Co(stage2_c26_c_fa1));
    FA fa_1007(.A(stage1_c25_c_fa6), .B(stage1_c25_c_fa7), .C(stage1_c25_c_ha0), .So(stage2_c26_s_fa2), .Co(stage2_c26_c_fa2));
    FA fa_1008(.A(stage1_c26_s_fa0), .B(stage1_c26_s_fa1), .C(stage1_c26_s_fa2), .So(stage2_c26_s_fa3), .Co(stage2_c26_c_fa3));
    FA fa_1009(.A(stage1_c26_s_fa3), .B(stage1_c26_s_fa4), .C(stage1_c26_s_fa5), .So(stage2_c26_s_fa4), .Co(stage2_c26_c_fa4));
    FA fa_1010(.A(stage1_c26_s_fa6), .B(stage1_c26_s_fa7), .C(stage1_c26_s_fa8), .So(stage2_c26_s_fa5), .Co(stage2_c26_c_fa5));
    FA fa_1011(.A(stage1_c26_c_fa0), .B(stage1_c26_c_fa1), .C(stage1_c26_c_fa2), .So(stage2_c27_s_fa0), .Co(stage2_c27_c_fa0));
    FA fa_1012(.A(stage1_c26_c_fa3), .B(stage1_c26_c_fa4), .C(stage1_c26_c_fa5), .So(stage2_c27_s_fa1), .Co(stage2_c27_c_fa1));
    FA fa_1013(.A(stage1_c26_c_fa6), .B(stage1_c26_c_fa7), .C(stage1_c26_c_fa8), .So(stage2_c27_s_fa2), .Co(stage2_c27_c_fa2));
    FA fa_1014(.A(stage1_c27_s_fa0), .B(stage1_c27_s_fa1), .C(stage1_c27_s_fa2), .So(stage2_c27_s_fa3), .Co(stage2_c27_c_fa3));
    FA fa_1015(.A(stage1_c27_s_fa3), .B(stage1_c27_s_fa4), .C(stage1_c27_s_fa5), .So(stage2_c27_s_fa4), .Co(stage2_c27_c_fa4));
    FA fa_1016(.A(stage1_c27_s_fa6), .B(stage1_c27_s_fa7), .C(stage1_c27_s_fa8), .So(stage2_c27_s_fa5), .Co(stage2_c27_c_fa5));
    FA fa_1017(.A(stage1_c27_c_fa0), .B(stage1_c27_c_fa1), .C(stage1_c27_c_fa2), .So(stage2_c28_s_fa0), .Co(stage2_c28_c_fa0));
    FA fa_1018(.A(stage1_c27_c_fa3), .B(stage1_c27_c_fa4), .C(stage1_c27_c_fa5), .So(stage2_c28_s_fa1), .Co(stage2_c28_c_fa1));
    FA fa_1019(.A(stage1_c27_c_fa6), .B(stage1_c27_c_fa7), .C(stage1_c27_c_fa8), .So(stage2_c28_s_fa2), .Co(stage2_c28_c_fa2));
    FA fa_1020(.A(stage1_c28_s_fa0), .B(stage1_c28_s_fa1), .C(stage1_c28_s_fa2), .So(stage2_c28_s_fa3), .Co(stage2_c28_c_fa3));
    FA fa_1021(.A(stage1_c28_s_fa3), .B(stage1_c28_s_fa4), .C(stage1_c28_s_fa5), .So(stage2_c28_s_fa4), .Co(stage2_c28_c_fa4));
    FA fa_1022(.A(stage1_c28_s_fa6), .B(stage1_c28_s_fa7), .C(stage1_c28_s_fa8), .So(stage2_c28_s_fa5), .Co(stage2_c28_c_fa5));
    FA fa_1023(.A(stage1_c28_c_fa0), .B(stage1_c28_c_fa1), .C(stage1_c28_c_fa2), .So(stage2_c29_s_fa0), .Co(stage2_c29_c_fa0));
    FA fa_1024(.A(stage1_c28_c_fa3), .B(stage1_c28_c_fa4), .C(stage1_c28_c_fa5), .So(stage2_c29_s_fa1), .Co(stage2_c29_c_fa1));
    FA fa_1025(.A(stage1_c28_c_fa6), .B(stage1_c28_c_fa7), .C(stage1_c28_c_fa8), .So(stage2_c29_s_fa2), .Co(stage2_c29_c_fa2));
    FA fa_1026(.A(stage1_c28_c_ha0), .B(stage1_c29_s_fa0), .C(stage1_c29_s_fa1), .So(stage2_c29_s_fa3), .Co(stage2_c29_c_fa3));
    FA fa_1027(.A(stage1_c29_s_fa2), .B(stage1_c29_s_fa3), .C(stage1_c29_s_fa4), .So(stage2_c29_s_fa4), .Co(stage2_c29_c_fa4));
    FA fa_1028(.A(stage1_c29_s_fa5), .B(stage1_c29_s_fa6), .C(stage1_c29_s_fa7), .So(stage2_c29_s_fa5), .Co(stage2_c29_c_fa5));
    HA ha_67(.A(stage1_c29_s_fa8), .B(stage1_c29_s_fa9), .So(stage2_c29_s_ha0), .Co(stage2_c29_c_ha0));
    FA fa_1029(.A(stage1_c29_c_fa0), .B(stage1_c29_c_fa1), .C(stage1_c29_c_fa2), .So(stage2_c30_s_fa0), .Co(stage2_c30_c_fa0));
    FA fa_1030(.A(stage1_c29_c_fa3), .B(stage1_c29_c_fa4), .C(stage1_c29_c_fa5), .So(stage2_c30_s_fa1), .Co(stage2_c30_c_fa1));
    FA fa_1031(.A(stage1_c29_c_fa6), .B(stage1_c29_c_fa7), .C(stage1_c29_c_fa8), .So(stage2_c30_s_fa2), .Co(stage2_c30_c_fa2));
    FA fa_1032(.A(stage1_c29_c_fa9), .B(stage1_c30_s_fa0), .C(stage1_c30_s_fa1), .So(stage2_c30_s_fa3), .Co(stage2_c30_c_fa3));
    FA fa_1033(.A(stage1_c30_s_fa2), .B(stage1_c30_s_fa3), .C(stage1_c30_s_fa4), .So(stage2_c30_s_fa4), .Co(stage2_c30_c_fa4));
    FA fa_1034(.A(stage1_c30_s_fa5), .B(stage1_c30_s_fa6), .C(stage1_c30_s_fa7), .So(stage2_c30_s_fa5), .Co(stage2_c30_c_fa5));
    FA fa_1035(.A(stage1_c30_s_fa8), .B(stage1_c30_s_fa9), .C(stage0_r30_c0), .So(stage2_c30_s_fa6), .Co(stage2_c30_c_fa6));
    FA fa_1036(.A(stage1_c30_c_fa0), .B(stage1_c30_c_fa1), .C(stage1_c30_c_fa2), .So(stage2_c31_s_fa0), .Co(stage2_c31_c_fa0));
    FA fa_1037(.A(stage1_c30_c_fa3), .B(stage1_c30_c_fa4), .C(stage1_c30_c_fa5), .So(stage2_c31_s_fa1), .Co(stage2_c31_c_fa1));
    FA fa_1038(.A(stage1_c30_c_fa6), .B(stage1_c30_c_fa7), .C(stage1_c30_c_fa8), .So(stage2_c31_s_fa2), .Co(stage2_c31_c_fa2));
    FA fa_1039(.A(stage1_c30_c_fa9), .B(stage1_c31_s_fa0), .C(stage1_c31_s_fa1), .So(stage2_c31_s_fa3), .Co(stage2_c31_c_fa3));
    FA fa_1040(.A(stage1_c31_s_fa2), .B(stage1_c31_s_fa3), .C(stage1_c31_s_fa4), .So(stage2_c31_s_fa4), .Co(stage2_c31_c_fa4));
    FA fa_1041(.A(stage1_c31_s_fa5), .B(stage1_c31_s_fa6), .C(stage1_c31_s_fa7), .So(stage2_c31_s_fa5), .Co(stage2_c31_c_fa5));
    FA fa_1042(.A(stage1_c31_s_fa8), .B(stage1_c31_s_fa9), .C(stage1_c31_s_ha0), .So(stage2_c31_s_fa6), .Co(stage2_c31_c_fa6));
    FA fa_1043(.A(stage1_c31_c_fa0), .B(stage1_c31_c_fa1), .C(stage1_c31_c_fa2), .So(stage2_c32_s_fa0), .Co(stage2_c32_c_fa0));
    FA fa_1044(.A(stage1_c31_c_fa3), .B(stage1_c31_c_fa4), .C(stage1_c31_c_fa5), .So(stage2_c32_s_fa1), .Co(stage2_c32_c_fa1));
    FA fa_1045(.A(stage1_c31_c_fa6), .B(stage1_c31_c_fa7), .C(stage1_c31_c_fa8), .So(stage2_c32_s_fa2), .Co(stage2_c32_c_fa2));
    FA fa_1046(.A(stage1_c31_c_fa9), .B(stage1_c31_c_ha0), .C(stage1_c32_s_fa0), .So(stage2_c32_s_fa3), .Co(stage2_c32_c_fa3));
    FA fa_1047(.A(stage1_c32_s_fa1), .B(stage1_c32_s_fa2), .C(stage1_c32_s_fa3), .So(stage2_c32_s_fa4), .Co(stage2_c32_c_fa4));
    FA fa_1048(.A(stage1_c32_s_fa4), .B(stage1_c32_s_fa5), .C(stage1_c32_s_fa6), .So(stage2_c32_s_fa5), .Co(stage2_c32_c_fa5));
    FA fa_1049(.A(stage1_c32_s_fa7), .B(stage1_c32_s_fa8), .C(stage1_c32_s_fa9), .So(stage2_c32_s_fa6), .Co(stage2_c32_c_fa6));
    FA fa_1050(.A(stage1_c32_c_fa0), .B(stage1_c32_c_fa1), .C(stage1_c32_c_fa2), .So(stage2_c33_s_fa0), .Co(stage2_c33_c_fa0));
    FA fa_1051(.A(stage1_c32_c_fa3), .B(stage1_c32_c_fa4), .C(stage1_c32_c_fa5), .So(stage2_c33_s_fa1), .Co(stage2_c33_c_fa1));
    FA fa_1052(.A(stage1_c32_c_fa6), .B(stage1_c32_c_fa7), .C(stage1_c32_c_fa8), .So(stage2_c33_s_fa2), .Co(stage2_c33_c_fa2));
    FA fa_1053(.A(stage1_c32_c_fa9), .B(stage1_c32_c_fa10), .C(stage1_c33_s_fa0), .So(stage2_c33_s_fa3), .Co(stage2_c33_c_fa3));
    FA fa_1054(.A(stage1_c33_s_fa1), .B(stage1_c33_s_fa2), .C(stage1_c33_s_fa3), .So(stage2_c33_s_fa4), .Co(stage2_c33_c_fa4));
    FA fa_1055(.A(stage1_c33_s_fa4), .B(stage1_c33_s_fa5), .C(stage1_c33_s_fa6), .So(stage2_c33_s_fa5), .Co(stage2_c33_c_fa5));
    FA fa_1056(.A(stage1_c33_s_fa7), .B(stage1_c33_s_fa8), .C(stage1_c33_s_fa9), .So(stage2_c33_s_fa6), .Co(stage2_c33_c_fa6));
    HA ha_68(.A(stage1_c33_s_fa10), .B(stage0_r33_c0), .So(stage2_c33_s_ha0), .Co(stage2_c33_c_ha0));
    FA fa_1057(.A(stage1_c33_c_fa0), .B(stage1_c33_c_fa1), .C(stage1_c33_c_fa2), .So(stage2_c34_s_fa0), .Co(stage2_c34_c_fa0));
    FA fa_1058(.A(stage1_c33_c_fa3), .B(stage1_c33_c_fa4), .C(stage1_c33_c_fa5), .So(stage2_c34_s_fa1), .Co(stage2_c34_c_fa1));
    FA fa_1059(.A(stage1_c33_c_fa6), .B(stage1_c33_c_fa7), .C(stage1_c33_c_fa8), .So(stage2_c34_s_fa2), .Co(stage2_c34_c_fa2));
    FA fa_1060(.A(stage1_c33_c_fa9), .B(stage1_c33_c_fa10), .C(stage1_c34_s_fa0), .So(stage2_c34_s_fa3), .Co(stage2_c34_c_fa3));
    FA fa_1061(.A(stage1_c34_s_fa1), .B(stage1_c34_s_fa2), .C(stage1_c34_s_fa3), .So(stage2_c34_s_fa4), .Co(stage2_c34_c_fa4));
    FA fa_1062(.A(stage1_c34_s_fa4), .B(stage1_c34_s_fa5), .C(stage1_c34_s_fa6), .So(stage2_c34_s_fa5), .Co(stage2_c34_c_fa5));
    FA fa_1063(.A(stage1_c34_s_fa7), .B(stage1_c34_s_fa8), .C(stage1_c34_s_fa9), .So(stage2_c34_s_fa6), .Co(stage2_c34_c_fa6));
    HA ha_69(.A(stage1_c34_s_fa10), .B(stage1_c34_s_ha0), .So(stage2_c34_s_ha0), .Co(stage2_c34_c_ha0));
    FA fa_1064(.A(stage1_c34_c_fa0), .B(stage1_c34_c_fa1), .C(stage1_c34_c_fa2), .So(stage2_c35_s_fa0), .Co(stage2_c35_c_fa0));
    FA fa_1065(.A(stage1_c34_c_fa3), .B(stage1_c34_c_fa4), .C(stage1_c34_c_fa5), .So(stage2_c35_s_fa1), .Co(stage2_c35_c_fa1));
    FA fa_1066(.A(stage1_c34_c_fa6), .B(stage1_c34_c_fa7), .C(stage1_c34_c_fa8), .So(stage2_c35_s_fa2), .Co(stage2_c35_c_fa2));
    FA fa_1067(.A(stage1_c34_c_fa9), .B(stage1_c34_c_fa10), .C(stage1_c34_c_ha0), .So(stage2_c35_s_fa3), .Co(stage2_c35_c_fa3));
    FA fa_1068(.A(stage1_c35_s_fa0), .B(stage1_c35_s_fa1), .C(stage1_c35_s_fa2), .So(stage2_c35_s_fa4), .Co(stage2_c35_c_fa4));
    FA fa_1069(.A(stage1_c35_s_fa3), .B(stage1_c35_s_fa4), .C(stage1_c35_s_fa5), .So(stage2_c35_s_fa5), .Co(stage2_c35_c_fa5));
    FA fa_1070(.A(stage1_c35_s_fa6), .B(stage1_c35_s_fa7), .C(stage1_c35_s_fa8), .So(stage2_c35_s_fa6), .Co(stage2_c35_c_fa6));
    FA fa_1071(.A(stage1_c35_s_fa9), .B(stage1_c35_s_fa10), .C(stage1_c35_s_fa11), .So(stage2_c35_s_fa7), .Co(stage2_c35_c_fa7));
    FA fa_1072(.A(stage1_c35_c_fa0), .B(stage1_c35_c_fa1), .C(stage1_c35_c_fa2), .So(stage2_c36_s_fa0), .Co(stage2_c36_c_fa0));
    FA fa_1073(.A(stage1_c35_c_fa3), .B(stage1_c35_c_fa4), .C(stage1_c35_c_fa5), .So(stage2_c36_s_fa1), .Co(stage2_c36_c_fa1));
    FA fa_1074(.A(stage1_c35_c_fa6), .B(stage1_c35_c_fa7), .C(stage1_c35_c_fa8), .So(stage2_c36_s_fa2), .Co(stage2_c36_c_fa2));
    FA fa_1075(.A(stage1_c35_c_fa9), .B(stage1_c35_c_fa10), .C(stage1_c35_c_fa11), .So(stage2_c36_s_fa3), .Co(stage2_c36_c_fa3));
    FA fa_1076(.A(stage1_c36_s_fa0), .B(stage1_c36_s_fa1), .C(stage1_c36_s_fa2), .So(stage2_c36_s_fa4), .Co(stage2_c36_c_fa4));
    FA fa_1077(.A(stage1_c36_s_fa3), .B(stage1_c36_s_fa4), .C(stage1_c36_s_fa5), .So(stage2_c36_s_fa5), .Co(stage2_c36_c_fa5));
    FA fa_1078(.A(stage1_c36_s_fa6), .B(stage1_c36_s_fa7), .C(stage1_c36_s_fa8), .So(stage2_c36_s_fa6), .Co(stage2_c36_c_fa6));
    FA fa_1079(.A(stage1_c36_s_fa9), .B(stage1_c36_s_fa10), .C(stage1_c36_s_fa11), .So(stage2_c36_s_fa7), .Co(stage2_c36_c_fa7));
    FA fa_1080(.A(stage1_c36_c_fa0), .B(stage1_c36_c_fa1), .C(stage1_c36_c_fa2), .So(stage2_c37_s_fa0), .Co(stage2_c37_c_fa0));
    FA fa_1081(.A(stage1_c36_c_fa3), .B(stage1_c36_c_fa4), .C(stage1_c36_c_fa5), .So(stage2_c37_s_fa1), .Co(stage2_c37_c_fa1));
    FA fa_1082(.A(stage1_c36_c_fa6), .B(stage1_c36_c_fa7), .C(stage1_c36_c_fa8), .So(stage2_c37_s_fa2), .Co(stage2_c37_c_fa2));
    FA fa_1083(.A(stage1_c36_c_fa9), .B(stage1_c36_c_fa10), .C(stage1_c36_c_fa11), .So(stage2_c37_s_fa3), .Co(stage2_c37_c_fa3));
    FA fa_1084(.A(stage1_c37_s_fa0), .B(stage1_c37_s_fa1), .C(stage1_c37_s_fa2), .So(stage2_c37_s_fa4), .Co(stage2_c37_c_fa4));
    FA fa_1085(.A(stage1_c37_s_fa3), .B(stage1_c37_s_fa4), .C(stage1_c37_s_fa5), .So(stage2_c37_s_fa5), .Co(stage2_c37_c_fa5));
    FA fa_1086(.A(stage1_c37_s_fa6), .B(stage1_c37_s_fa7), .C(stage1_c37_s_fa8), .So(stage2_c37_s_fa6), .Co(stage2_c37_c_fa6));
    FA fa_1087(.A(stage1_c37_s_fa9), .B(stage1_c37_s_fa10), .C(stage1_c37_s_fa11), .So(stage2_c37_s_fa7), .Co(stage2_c37_c_fa7));
    FA fa_1088(.A(stage1_c37_c_fa0), .B(stage1_c37_c_fa1), .C(stage1_c37_c_fa2), .So(stage2_c38_s_fa0), .Co(stage2_c38_c_fa0));
    FA fa_1089(.A(stage1_c37_c_fa3), .B(stage1_c37_c_fa4), .C(stage1_c37_c_fa5), .So(stage2_c38_s_fa1), .Co(stage2_c38_c_fa1));
    FA fa_1090(.A(stage1_c37_c_fa6), .B(stage1_c37_c_fa7), .C(stage1_c37_c_fa8), .So(stage2_c38_s_fa2), .Co(stage2_c38_c_fa2));
    FA fa_1091(.A(stage1_c37_c_fa9), .B(stage1_c37_c_fa10), .C(stage1_c37_c_fa11), .So(stage2_c38_s_fa3), .Co(stage2_c38_c_fa3));
    FA fa_1092(.A(stage1_c37_c_ha0), .B(stage1_c38_s_fa0), .C(stage1_c38_s_fa1), .So(stage2_c38_s_fa4), .Co(stage2_c38_c_fa4));
    FA fa_1093(.A(stage1_c38_s_fa2), .B(stage1_c38_s_fa3), .C(stage1_c38_s_fa4), .So(stage2_c38_s_fa5), .Co(stage2_c38_c_fa5));
    FA fa_1094(.A(stage1_c38_s_fa5), .B(stage1_c38_s_fa6), .C(stage1_c38_s_fa7), .So(stage2_c38_s_fa6), .Co(stage2_c38_c_fa6));
    FA fa_1095(.A(stage1_c38_s_fa8), .B(stage1_c38_s_fa9), .C(stage1_c38_s_fa10), .So(stage2_c38_s_fa7), .Co(stage2_c38_c_fa7));
    HA ha_70(.A(stage1_c38_s_fa11), .B(stage1_c38_s_fa12), .So(stage2_c38_s_ha0), .Co(stage2_c38_c_ha0));
    FA fa_1096(.A(stage1_c38_c_fa0), .B(stage1_c38_c_fa1), .C(stage1_c38_c_fa2), .So(stage2_c39_s_fa0), .Co(stage2_c39_c_fa0));
    FA fa_1097(.A(stage1_c38_c_fa3), .B(stage1_c38_c_fa4), .C(stage1_c38_c_fa5), .So(stage2_c39_s_fa1), .Co(stage2_c39_c_fa1));
    FA fa_1098(.A(stage1_c38_c_fa6), .B(stage1_c38_c_fa7), .C(stage1_c38_c_fa8), .So(stage2_c39_s_fa2), .Co(stage2_c39_c_fa2));
    FA fa_1099(.A(stage1_c38_c_fa9), .B(stage1_c38_c_fa10), .C(stage1_c38_c_fa11), .So(stage2_c39_s_fa3), .Co(stage2_c39_c_fa3));
    FA fa_1100(.A(stage1_c38_c_fa12), .B(stage1_c39_s_fa0), .C(stage1_c39_s_fa1), .So(stage2_c39_s_fa4), .Co(stage2_c39_c_fa4));
    FA fa_1101(.A(stage1_c39_s_fa2), .B(stage1_c39_s_fa3), .C(stage1_c39_s_fa4), .So(stage2_c39_s_fa5), .Co(stage2_c39_c_fa5));
    FA fa_1102(.A(stage1_c39_s_fa5), .B(stage1_c39_s_fa6), .C(stage1_c39_s_fa7), .So(stage2_c39_s_fa6), .Co(stage2_c39_c_fa6));
    FA fa_1103(.A(stage1_c39_s_fa8), .B(stage1_c39_s_fa9), .C(stage1_c39_s_fa10), .So(stage2_c39_s_fa7), .Co(stage2_c39_c_fa7));
    FA fa_1104(.A(stage1_c39_s_fa11), .B(stage1_c39_s_fa12), .C(stage0_r39_c0), .So(stage2_c39_s_fa8), .Co(stage2_c39_c_fa8));
    FA fa_1105(.A(stage1_c39_c_fa0), .B(stage1_c39_c_fa1), .C(stage1_c39_c_fa2), .So(stage2_c40_s_fa0), .Co(stage2_c40_c_fa0));
    FA fa_1106(.A(stage1_c39_c_fa3), .B(stage1_c39_c_fa4), .C(stage1_c39_c_fa5), .So(stage2_c40_s_fa1), .Co(stage2_c40_c_fa1));
    FA fa_1107(.A(stage1_c39_c_fa6), .B(stage1_c39_c_fa7), .C(stage1_c39_c_fa8), .So(stage2_c40_s_fa2), .Co(stage2_c40_c_fa2));
    FA fa_1108(.A(stage1_c39_c_fa9), .B(stage1_c39_c_fa10), .C(stage1_c39_c_fa11), .So(stage2_c40_s_fa3), .Co(stage2_c40_c_fa3));
    FA fa_1109(.A(stage1_c39_c_fa12), .B(stage1_c40_s_fa0), .C(stage1_c40_s_fa1), .So(stage2_c40_s_fa4), .Co(stage2_c40_c_fa4));
    FA fa_1110(.A(stage1_c40_s_fa2), .B(stage1_c40_s_fa3), .C(stage1_c40_s_fa4), .So(stage2_c40_s_fa5), .Co(stage2_c40_c_fa5));
    FA fa_1111(.A(stage1_c40_s_fa5), .B(stage1_c40_s_fa6), .C(stage1_c40_s_fa7), .So(stage2_c40_s_fa6), .Co(stage2_c40_c_fa6));
    FA fa_1112(.A(stage1_c40_s_fa8), .B(stage1_c40_s_fa9), .C(stage1_c40_s_fa10), .So(stage2_c40_s_fa7), .Co(stage2_c40_c_fa7));
    FA fa_1113(.A(stage1_c40_s_fa11), .B(stage1_c40_s_fa12), .C(stage1_c40_s_ha0), .So(stage2_c40_s_fa8), .Co(stage2_c40_c_fa8));
    FA fa_1114(.A(stage1_c40_c_fa0), .B(stage1_c40_c_fa1), .C(stage1_c40_c_fa2), .So(stage2_c41_s_fa0), .Co(stage2_c41_c_fa0));
    FA fa_1115(.A(stage1_c40_c_fa3), .B(stage1_c40_c_fa4), .C(stage1_c40_c_fa5), .So(stage2_c41_s_fa1), .Co(stage2_c41_c_fa1));
    FA fa_1116(.A(stage1_c40_c_fa6), .B(stage1_c40_c_fa7), .C(stage1_c40_c_fa8), .So(stage2_c41_s_fa2), .Co(stage2_c41_c_fa2));
    FA fa_1117(.A(stage1_c40_c_fa9), .B(stage1_c40_c_fa10), .C(stage1_c40_c_fa11), .So(stage2_c41_s_fa3), .Co(stage2_c41_c_fa3));
    FA fa_1118(.A(stage1_c40_c_fa12), .B(stage1_c40_c_ha0), .C(stage1_c41_s_fa0), .So(stage2_c41_s_fa4), .Co(stage2_c41_c_fa4));
    FA fa_1119(.A(stage1_c41_s_fa1), .B(stage1_c41_s_fa2), .C(stage1_c41_s_fa3), .So(stage2_c41_s_fa5), .Co(stage2_c41_c_fa5));
    FA fa_1120(.A(stage1_c41_s_fa4), .B(stage1_c41_s_fa5), .C(stage1_c41_s_fa6), .So(stage2_c41_s_fa6), .Co(stage2_c41_c_fa6));
    FA fa_1121(.A(stage1_c41_s_fa7), .B(stage1_c41_s_fa8), .C(stage1_c41_s_fa9), .So(stage2_c41_s_fa7), .Co(stage2_c41_c_fa7));
    FA fa_1122(.A(stage1_c41_s_fa10), .B(stage1_c41_s_fa11), .C(stage1_c41_s_fa12), .So(stage2_c41_s_fa8), .Co(stage2_c41_c_fa8));
    FA fa_1123(.A(stage1_c41_c_fa0), .B(stage1_c41_c_fa1), .C(stage1_c41_c_fa2), .So(stage2_c42_s_fa0), .Co(stage2_c42_c_fa0));
    FA fa_1124(.A(stage1_c41_c_fa3), .B(stage1_c41_c_fa4), .C(stage1_c41_c_fa5), .So(stage2_c42_s_fa1), .Co(stage2_c42_c_fa1));
    FA fa_1125(.A(stage1_c41_c_fa6), .B(stage1_c41_c_fa7), .C(stage1_c41_c_fa8), .So(stage2_c42_s_fa2), .Co(stage2_c42_c_fa2));
    FA fa_1126(.A(stage1_c41_c_fa9), .B(stage1_c41_c_fa10), .C(stage1_c41_c_fa11), .So(stage2_c42_s_fa3), .Co(stage2_c42_c_fa3));
    FA fa_1127(.A(stage1_c41_c_fa12), .B(stage1_c41_c_ha0), .C(stage1_c42_s_fa0), .So(stage2_c42_s_fa4), .Co(stage2_c42_c_fa4));
    FA fa_1128(.A(stage1_c42_s_fa1), .B(stage1_c42_s_fa2), .C(stage1_c42_s_fa3), .So(stage2_c42_s_fa5), .Co(stage2_c42_c_fa5));
    FA fa_1129(.A(stage1_c42_s_fa4), .B(stage1_c42_s_fa5), .C(stage1_c42_s_fa6), .So(stage2_c42_s_fa6), .Co(stage2_c42_c_fa6));
    FA fa_1130(.A(stage1_c42_s_fa7), .B(stage1_c42_s_fa8), .C(stage1_c42_s_fa9), .So(stage2_c42_s_fa7), .Co(stage2_c42_c_fa7));
    FA fa_1131(.A(stage1_c42_s_fa10), .B(stage1_c42_s_fa11), .C(stage1_c42_s_fa12), .So(stage2_c42_s_fa8), .Co(stage2_c42_c_fa8));
    FA fa_1132(.A(stage1_c42_c_fa0), .B(stage1_c42_c_fa1), .C(stage1_c42_c_fa2), .So(stage2_c43_s_fa0), .Co(stage2_c43_c_fa0));
    FA fa_1133(.A(stage1_c42_c_fa3), .B(stage1_c42_c_fa4), .C(stage1_c42_c_fa5), .So(stage2_c43_s_fa1), .Co(stage2_c43_c_fa1));
    FA fa_1134(.A(stage1_c42_c_fa6), .B(stage1_c42_c_fa7), .C(stage1_c42_c_fa8), .So(stage2_c43_s_fa2), .Co(stage2_c43_c_fa2));
    FA fa_1135(.A(stage1_c42_c_fa9), .B(stage1_c42_c_fa10), .C(stage1_c42_c_fa11), .So(stage2_c43_s_fa3), .Co(stage2_c43_c_fa3));
    FA fa_1136(.A(stage1_c42_c_fa12), .B(stage1_c42_c_ha0), .C(stage1_c43_s_fa0), .So(stage2_c43_s_fa4), .Co(stage2_c43_c_fa4));
    FA fa_1137(.A(stage1_c43_s_fa1), .B(stage1_c43_s_fa2), .C(stage1_c43_s_fa3), .So(stage2_c43_s_fa5), .Co(stage2_c43_c_fa5));
    FA fa_1138(.A(stage1_c43_s_fa4), .B(stage1_c43_s_fa5), .C(stage1_c43_s_fa6), .So(stage2_c43_s_fa6), .Co(stage2_c43_c_fa6));
    FA fa_1139(.A(stage1_c43_s_fa7), .B(stage1_c43_s_fa8), .C(stage1_c43_s_fa9), .So(stage2_c43_s_fa7), .Co(stage2_c43_c_fa7));
    FA fa_1140(.A(stage1_c43_s_fa10), .B(stage1_c43_s_fa11), .C(stage1_c43_s_fa12), .So(stage2_c43_s_fa8), .Co(stage2_c43_c_fa8));
    FA fa_1141(.A(stage1_c43_c_fa0), .B(stage1_c43_c_fa1), .C(stage1_c43_c_fa2), .So(stage2_c44_s_fa0), .Co(stage2_c44_c_fa0));
    FA fa_1142(.A(stage1_c43_c_fa3), .B(stage1_c43_c_fa4), .C(stage1_c43_c_fa5), .So(stage2_c44_s_fa1), .Co(stage2_c44_c_fa1));
    FA fa_1143(.A(stage1_c43_c_fa6), .B(stage1_c43_c_fa7), .C(stage1_c43_c_fa8), .So(stage2_c44_s_fa2), .Co(stage2_c44_c_fa2));
    FA fa_1144(.A(stage1_c43_c_fa9), .B(stage1_c43_c_fa10), .C(stage1_c43_c_fa11), .So(stage2_c44_s_fa3), .Co(stage2_c44_c_fa3));
    FA fa_1145(.A(stage1_c43_c_fa12), .B(stage1_c43_c_ha0), .C(stage1_c44_s_fa0), .So(stage2_c44_s_fa4), .Co(stage2_c44_c_fa4));
    FA fa_1146(.A(stage1_c44_s_fa1), .B(stage1_c44_s_fa2), .C(stage1_c44_s_fa3), .So(stage2_c44_s_fa5), .Co(stage2_c44_c_fa5));
    FA fa_1147(.A(stage1_c44_s_fa4), .B(stage1_c44_s_fa5), .C(stage1_c44_s_fa6), .So(stage2_c44_s_fa6), .Co(stage2_c44_c_fa6));
    FA fa_1148(.A(stage1_c44_s_fa7), .B(stage1_c44_s_fa8), .C(stage1_c44_s_fa9), .So(stage2_c44_s_fa7), .Co(stage2_c44_c_fa7));
    FA fa_1149(.A(stage1_c44_s_fa10), .B(stage1_c44_s_fa11), .C(stage1_c44_s_fa12), .So(stage2_c44_s_fa8), .Co(stage2_c44_c_fa8));
    FA fa_1150(.A(stage1_c44_c_fa0), .B(stage1_c44_c_fa1), .C(stage1_c44_c_fa2), .So(stage2_c45_s_fa0), .Co(stage2_c45_c_fa0));
    FA fa_1151(.A(stage1_c44_c_fa3), .B(stage1_c44_c_fa4), .C(stage1_c44_c_fa5), .So(stage2_c45_s_fa1), .Co(stage2_c45_c_fa1));
    FA fa_1152(.A(stage1_c44_c_fa6), .B(stage1_c44_c_fa7), .C(stage1_c44_c_fa8), .So(stage2_c45_s_fa2), .Co(stage2_c45_c_fa2));
    FA fa_1153(.A(stage1_c44_c_fa9), .B(stage1_c44_c_fa10), .C(stage1_c44_c_fa11), .So(stage2_c45_s_fa3), .Co(stage2_c45_c_fa3));
    FA fa_1154(.A(stage1_c44_c_fa12), .B(stage1_c44_c_ha0), .C(stage1_c45_s_fa0), .So(stage2_c45_s_fa4), .Co(stage2_c45_c_fa4));
    FA fa_1155(.A(stage1_c45_s_fa1), .B(stage1_c45_s_fa2), .C(stage1_c45_s_fa3), .So(stage2_c45_s_fa5), .Co(stage2_c45_c_fa5));
    FA fa_1156(.A(stage1_c45_s_fa4), .B(stage1_c45_s_fa5), .C(stage1_c45_s_fa6), .So(stage2_c45_s_fa6), .Co(stage2_c45_c_fa6));
    FA fa_1157(.A(stage1_c45_s_fa7), .B(stage1_c45_s_fa8), .C(stage1_c45_s_fa9), .So(stage2_c45_s_fa7), .Co(stage2_c45_c_fa7));
    FA fa_1158(.A(stage1_c45_s_fa10), .B(stage1_c45_s_fa11), .C(stage1_c45_s_fa12), .So(stage2_c45_s_fa8), .Co(stage2_c45_c_fa8));
    FA fa_1159(.A(stage1_c45_c_fa0), .B(stage1_c45_c_fa1), .C(stage1_c45_c_fa2), .So(stage2_c46_s_fa0), .Co(stage2_c46_c_fa0));
    FA fa_1160(.A(stage1_c45_c_fa3), .B(stage1_c45_c_fa4), .C(stage1_c45_c_fa5), .So(stage2_c46_s_fa1), .Co(stage2_c46_c_fa1));
    FA fa_1161(.A(stage1_c45_c_fa6), .B(stage1_c45_c_fa7), .C(stage1_c45_c_fa8), .So(stage2_c46_s_fa2), .Co(stage2_c46_c_fa2));
    FA fa_1162(.A(stage1_c45_c_fa9), .B(stage1_c45_c_fa10), .C(stage1_c45_c_fa11), .So(stage2_c46_s_fa3), .Co(stage2_c46_c_fa3));
    FA fa_1163(.A(stage1_c45_c_fa12), .B(stage1_c45_c_ha0), .C(stage1_c46_s_fa0), .So(stage2_c46_s_fa4), .Co(stage2_c46_c_fa4));
    FA fa_1164(.A(stage1_c46_s_fa1), .B(stage1_c46_s_fa2), .C(stage1_c46_s_fa3), .So(stage2_c46_s_fa5), .Co(stage2_c46_c_fa5));
    FA fa_1165(.A(stage1_c46_s_fa4), .B(stage1_c46_s_fa5), .C(stage1_c46_s_fa6), .So(stage2_c46_s_fa6), .Co(stage2_c46_c_fa6));
    FA fa_1166(.A(stage1_c46_s_fa7), .B(stage1_c46_s_fa8), .C(stage1_c46_s_fa9), .So(stage2_c46_s_fa7), .Co(stage2_c46_c_fa7));
    FA fa_1167(.A(stage1_c46_s_fa10), .B(stage1_c46_s_fa11), .C(stage1_c46_s_fa12), .So(stage2_c46_s_fa8), .Co(stage2_c46_c_fa8));
    FA fa_1168(.A(stage1_c46_c_fa0), .B(stage1_c46_c_fa1), .C(stage1_c46_c_fa2), .So(stage2_c47_s_fa0), .Co(stage2_c47_c_fa0));
    FA fa_1169(.A(stage1_c46_c_fa3), .B(stage1_c46_c_fa4), .C(stage1_c46_c_fa5), .So(stage2_c47_s_fa1), .Co(stage2_c47_c_fa1));
    FA fa_1170(.A(stage1_c46_c_fa6), .B(stage1_c46_c_fa7), .C(stage1_c46_c_fa8), .So(stage2_c47_s_fa2), .Co(stage2_c47_c_fa2));
    FA fa_1171(.A(stage1_c46_c_fa9), .B(stage1_c46_c_fa10), .C(stage1_c46_c_fa11), .So(stage2_c47_s_fa3), .Co(stage2_c47_c_fa3));
    FA fa_1172(.A(stage1_c46_c_fa12), .B(stage1_c46_c_ha0), .C(stage1_c47_s_fa0), .So(stage2_c47_s_fa4), .Co(stage2_c47_c_fa4));
    FA fa_1173(.A(stage1_c47_s_fa1), .B(stage1_c47_s_fa2), .C(stage1_c47_s_fa3), .So(stage2_c47_s_fa5), .Co(stage2_c47_c_fa5));
    FA fa_1174(.A(stage1_c47_s_fa4), .B(stage1_c47_s_fa5), .C(stage1_c47_s_fa6), .So(stage2_c47_s_fa6), .Co(stage2_c47_c_fa6));
    FA fa_1175(.A(stage1_c47_s_fa7), .B(stage1_c47_s_fa8), .C(stage1_c47_s_fa9), .So(stage2_c47_s_fa7), .Co(stage2_c47_c_fa7));
    FA fa_1176(.A(stage1_c47_s_fa10), .B(stage1_c47_s_fa11), .C(stage1_c47_s_fa12), .So(stage2_c47_s_fa8), .Co(stage2_c47_c_fa8));
    FA fa_1177(.A(stage1_c47_c_fa0), .B(stage1_c47_c_fa1), .C(stage1_c47_c_fa2), .So(stage2_c48_s_fa0), .Co(stage2_c48_c_fa0));
    FA fa_1178(.A(stage1_c47_c_fa3), .B(stage1_c47_c_fa4), .C(stage1_c47_c_fa5), .So(stage2_c48_s_fa1), .Co(stage2_c48_c_fa1));
    FA fa_1179(.A(stage1_c47_c_fa6), .B(stage1_c47_c_fa7), .C(stage1_c47_c_fa8), .So(stage2_c48_s_fa2), .Co(stage2_c48_c_fa2));
    FA fa_1180(.A(stage1_c47_c_fa9), .B(stage1_c47_c_fa10), .C(stage1_c47_c_fa11), .So(stage2_c48_s_fa3), .Co(stage2_c48_c_fa3));
    FA fa_1181(.A(stage1_c47_c_fa12), .B(stage1_c47_c_ha0), .C(stage1_c48_s_fa0), .So(stage2_c48_s_fa4), .Co(stage2_c48_c_fa4));
    FA fa_1182(.A(stage1_c48_s_fa1), .B(stage1_c48_s_fa2), .C(stage1_c48_s_fa3), .So(stage2_c48_s_fa5), .Co(stage2_c48_c_fa5));
    FA fa_1183(.A(stage1_c48_s_fa4), .B(stage1_c48_s_fa5), .C(stage1_c48_s_fa6), .So(stage2_c48_s_fa6), .Co(stage2_c48_c_fa6));
    FA fa_1184(.A(stage1_c48_s_fa7), .B(stage1_c48_s_fa8), .C(stage1_c48_s_fa9), .So(stage2_c48_s_fa7), .Co(stage2_c48_c_fa7));
    FA fa_1185(.A(stage1_c48_s_fa10), .B(stage1_c48_s_fa11), .C(stage1_c48_s_fa12), .So(stage2_c48_s_fa8), .Co(stage2_c48_c_fa8));
    FA fa_1186(.A(stage1_c48_c_fa0), .B(stage1_c48_c_fa1), .C(stage1_c48_c_fa2), .So(stage2_c49_s_fa0), .Co(stage2_c49_c_fa0));
    FA fa_1187(.A(stage1_c48_c_fa3), .B(stage1_c48_c_fa4), .C(stage1_c48_c_fa5), .So(stage2_c49_s_fa1), .Co(stage2_c49_c_fa1));
    FA fa_1188(.A(stage1_c48_c_fa6), .B(stage1_c48_c_fa7), .C(stage1_c48_c_fa8), .So(stage2_c49_s_fa2), .Co(stage2_c49_c_fa2));
    FA fa_1189(.A(stage1_c48_c_fa9), .B(stage1_c48_c_fa10), .C(stage1_c48_c_fa11), .So(stage2_c49_s_fa3), .Co(stage2_c49_c_fa3));
    FA fa_1190(.A(stage1_c48_c_fa12), .B(stage1_c48_c_ha0), .C(stage1_c49_s_fa0), .So(stage2_c49_s_fa4), .Co(stage2_c49_c_fa4));
    FA fa_1191(.A(stage1_c49_s_fa1), .B(stage1_c49_s_fa2), .C(stage1_c49_s_fa3), .So(stage2_c49_s_fa5), .Co(stage2_c49_c_fa5));
    FA fa_1192(.A(stage1_c49_s_fa4), .B(stage1_c49_s_fa5), .C(stage1_c49_s_fa6), .So(stage2_c49_s_fa6), .Co(stage2_c49_c_fa6));
    FA fa_1193(.A(stage1_c49_s_fa7), .B(stage1_c49_s_fa8), .C(stage1_c49_s_fa9), .So(stage2_c49_s_fa7), .Co(stage2_c49_c_fa7));
    FA fa_1194(.A(stage1_c49_s_fa10), .B(stage1_c49_s_fa11), .C(stage1_c49_s_fa12), .So(stage2_c49_s_fa8), .Co(stage2_c49_c_fa8));
    FA fa_1195(.A(stage1_c49_c_fa0), .B(stage1_c49_c_fa1), .C(stage1_c49_c_fa2), .So(stage2_c50_s_fa0), .Co(stage2_c50_c_fa0));
    FA fa_1196(.A(stage1_c49_c_fa3), .B(stage1_c49_c_fa4), .C(stage1_c49_c_fa5), .So(stage2_c50_s_fa1), .Co(stage2_c50_c_fa1));
    FA fa_1197(.A(stage1_c49_c_fa6), .B(stage1_c49_c_fa7), .C(stage1_c49_c_fa8), .So(stage2_c50_s_fa2), .Co(stage2_c50_c_fa2));
    FA fa_1198(.A(stage1_c49_c_fa9), .B(stage1_c49_c_fa10), .C(stage1_c49_c_fa11), .So(stage2_c50_s_fa3), .Co(stage2_c50_c_fa3));
    FA fa_1199(.A(stage1_c49_c_fa12), .B(stage1_c49_c_ha0), .C(stage1_c50_s_fa0), .So(stage2_c50_s_fa4), .Co(stage2_c50_c_fa4));
    FA fa_1200(.A(stage1_c50_s_fa1), .B(stage1_c50_s_fa2), .C(stage1_c50_s_fa3), .So(stage2_c50_s_fa5), .Co(stage2_c50_c_fa5));
    FA fa_1201(.A(stage1_c50_s_fa4), .B(stage1_c50_s_fa5), .C(stage1_c50_s_fa6), .So(stage2_c50_s_fa6), .Co(stage2_c50_c_fa6));
    FA fa_1202(.A(stage1_c50_s_fa7), .B(stage1_c50_s_fa8), .C(stage1_c50_s_fa9), .So(stage2_c50_s_fa7), .Co(stage2_c50_c_fa7));
    FA fa_1203(.A(stage1_c50_s_fa10), .B(stage1_c50_s_fa11), .C(stage1_c50_s_fa12), .So(stage2_c50_s_fa8), .Co(stage2_c50_c_fa8));
    FA fa_1204(.A(stage1_c50_c_fa0), .B(stage1_c50_c_fa1), .C(stage1_c50_c_fa2), .So(stage2_c51_s_fa0), .Co(stage2_c51_c_fa0));
    FA fa_1205(.A(stage1_c50_c_fa3), .B(stage1_c50_c_fa4), .C(stage1_c50_c_fa5), .So(stage2_c51_s_fa1), .Co(stage2_c51_c_fa1));
    FA fa_1206(.A(stage1_c50_c_fa6), .B(stage1_c50_c_fa7), .C(stage1_c50_c_fa8), .So(stage2_c51_s_fa2), .Co(stage2_c51_c_fa2));
    FA fa_1207(.A(stage1_c50_c_fa9), .B(stage1_c50_c_fa10), .C(stage1_c50_c_fa11), .So(stage2_c51_s_fa3), .Co(stage2_c51_c_fa3));
    FA fa_1208(.A(stage1_c50_c_fa12), .B(stage1_c50_c_ha0), .C(stage1_c51_s_fa0), .So(stage2_c51_s_fa4), .Co(stage2_c51_c_fa4));
    FA fa_1209(.A(stage1_c51_s_fa1), .B(stage1_c51_s_fa2), .C(stage1_c51_s_fa3), .So(stage2_c51_s_fa5), .Co(stage2_c51_c_fa5));
    FA fa_1210(.A(stage1_c51_s_fa4), .B(stage1_c51_s_fa5), .C(stage1_c51_s_fa6), .So(stage2_c51_s_fa6), .Co(stage2_c51_c_fa6));
    FA fa_1211(.A(stage1_c51_s_fa7), .B(stage1_c51_s_fa8), .C(stage1_c51_s_fa9), .So(stage2_c51_s_fa7), .Co(stage2_c51_c_fa7));
    FA fa_1212(.A(stage1_c51_s_fa10), .B(stage1_c51_s_fa11), .C(stage1_c51_s_fa12), .So(stage2_c51_s_fa8), .Co(stage2_c51_c_fa8));
    FA fa_1213(.A(stage1_c51_c_fa0), .B(stage1_c51_c_fa1), .C(stage1_c51_c_fa2), .So(stage2_c52_s_fa0), .Co(stage2_c52_c_fa0));
    FA fa_1214(.A(stage1_c51_c_fa3), .B(stage1_c51_c_fa4), .C(stage1_c51_c_fa5), .So(stage2_c52_s_fa1), .Co(stage2_c52_c_fa1));
    FA fa_1215(.A(stage1_c51_c_fa6), .B(stage1_c51_c_fa7), .C(stage1_c51_c_fa8), .So(stage2_c52_s_fa2), .Co(stage2_c52_c_fa2));
    FA fa_1216(.A(stage1_c51_c_fa9), .B(stage1_c51_c_fa10), .C(stage1_c51_c_fa11), .So(stage2_c52_s_fa3), .Co(stage2_c52_c_fa3));
    FA fa_1217(.A(stage1_c51_c_fa12), .B(stage1_c51_c_ha0), .C(stage1_c52_s_fa0), .So(stage2_c52_s_fa4), .Co(stage2_c52_c_fa4));
    FA fa_1218(.A(stage1_c52_s_fa1), .B(stage1_c52_s_fa2), .C(stage1_c52_s_fa3), .So(stage2_c52_s_fa5), .Co(stage2_c52_c_fa5));
    FA fa_1219(.A(stage1_c52_s_fa4), .B(stage1_c52_s_fa5), .C(stage1_c52_s_fa6), .So(stage2_c52_s_fa6), .Co(stage2_c52_c_fa6));
    FA fa_1220(.A(stage1_c52_s_fa7), .B(stage1_c52_s_fa8), .C(stage1_c52_s_fa9), .So(stage2_c52_s_fa7), .Co(stage2_c52_c_fa7));
    FA fa_1221(.A(stage1_c52_s_fa10), .B(stage1_c52_s_fa11), .C(stage1_c52_s_fa12), .So(stage2_c52_s_fa8), .Co(stage2_c52_c_fa8));
    FA fa_1222(.A(stage1_c52_c_fa0), .B(stage1_c52_c_fa1), .C(stage1_c52_c_fa2), .So(stage2_c53_s_fa0), .Co(stage2_c53_c_fa0));
    FA fa_1223(.A(stage1_c52_c_fa3), .B(stage1_c52_c_fa4), .C(stage1_c52_c_fa5), .So(stage2_c53_s_fa1), .Co(stage2_c53_c_fa1));
    FA fa_1224(.A(stage1_c52_c_fa6), .B(stage1_c52_c_fa7), .C(stage1_c52_c_fa8), .So(stage2_c53_s_fa2), .Co(stage2_c53_c_fa2));
    FA fa_1225(.A(stage1_c52_c_fa9), .B(stage1_c52_c_fa10), .C(stage1_c52_c_fa11), .So(stage2_c53_s_fa3), .Co(stage2_c53_c_fa3));
    FA fa_1226(.A(stage1_c52_c_fa12), .B(stage1_c52_c_ha0), .C(stage1_c53_s_fa0), .So(stage2_c53_s_fa4), .Co(stage2_c53_c_fa4));
    FA fa_1227(.A(stage1_c53_s_fa1), .B(stage1_c53_s_fa2), .C(stage1_c53_s_fa3), .So(stage2_c53_s_fa5), .Co(stage2_c53_c_fa5));
    FA fa_1228(.A(stage1_c53_s_fa4), .B(stage1_c53_s_fa5), .C(stage1_c53_s_fa6), .So(stage2_c53_s_fa6), .Co(stage2_c53_c_fa6));
    FA fa_1229(.A(stage1_c53_s_fa7), .B(stage1_c53_s_fa8), .C(stage1_c53_s_fa9), .So(stage2_c53_s_fa7), .Co(stage2_c53_c_fa7));
    FA fa_1230(.A(stage1_c53_s_fa10), .B(stage1_c53_s_fa11), .C(stage1_c53_s_fa12), .So(stage2_c53_s_fa8), .Co(stage2_c53_c_fa8));
    FA fa_1231(.A(stage1_c53_c_fa0), .B(stage1_c53_c_fa1), .C(stage1_c53_c_fa2), .So(stage2_c54_s_fa0), .Co(stage2_c54_c_fa0));
    FA fa_1232(.A(stage1_c53_c_fa3), .B(stage1_c53_c_fa4), .C(stage1_c53_c_fa5), .So(stage2_c54_s_fa1), .Co(stage2_c54_c_fa1));
    FA fa_1233(.A(stage1_c53_c_fa6), .B(stage1_c53_c_fa7), .C(stage1_c53_c_fa8), .So(stage2_c54_s_fa2), .Co(stage2_c54_c_fa2));
    FA fa_1234(.A(stage1_c53_c_fa9), .B(stage1_c53_c_fa10), .C(stage1_c53_c_fa11), .So(stage2_c54_s_fa3), .Co(stage2_c54_c_fa3));
    FA fa_1235(.A(stage1_c53_c_fa12), .B(stage1_c53_c_ha0), .C(stage1_c54_s_fa0), .So(stage2_c54_s_fa4), .Co(stage2_c54_c_fa4));
    FA fa_1236(.A(stage1_c54_s_fa1), .B(stage1_c54_s_fa2), .C(stage1_c54_s_fa3), .So(stage2_c54_s_fa5), .Co(stage2_c54_c_fa5));
    FA fa_1237(.A(stage1_c54_s_fa4), .B(stage1_c54_s_fa5), .C(stage1_c54_s_fa6), .So(stage2_c54_s_fa6), .Co(stage2_c54_c_fa6));
    FA fa_1238(.A(stage1_c54_s_fa7), .B(stage1_c54_s_fa8), .C(stage1_c54_s_fa9), .So(stage2_c54_s_fa7), .Co(stage2_c54_c_fa7));
    FA fa_1239(.A(stage1_c54_s_fa10), .B(stage1_c54_s_fa11), .C(stage1_c54_s_fa12), .So(stage2_c54_s_fa8), .Co(stage2_c54_c_fa8));
    FA fa_1240(.A(stage1_c54_c_fa0), .B(stage1_c54_c_fa1), .C(stage1_c54_c_fa2), .So(stage2_c55_s_fa0), .Co(stage2_c55_c_fa0));
    FA fa_1241(.A(stage1_c54_c_fa3), .B(stage1_c54_c_fa4), .C(stage1_c54_c_fa5), .So(stage2_c55_s_fa1), .Co(stage2_c55_c_fa1));
    FA fa_1242(.A(stage1_c54_c_fa6), .B(stage1_c54_c_fa7), .C(stage1_c54_c_fa8), .So(stage2_c55_s_fa2), .Co(stage2_c55_c_fa2));
    FA fa_1243(.A(stage1_c54_c_fa9), .B(stage1_c54_c_fa10), .C(stage1_c54_c_fa11), .So(stage2_c55_s_fa3), .Co(stage2_c55_c_fa3));
    FA fa_1244(.A(stage1_c54_c_fa12), .B(stage1_c54_c_ha0), .C(stage1_c55_s_fa0), .So(stage2_c55_s_fa4), .Co(stage2_c55_c_fa4));
    FA fa_1245(.A(stage1_c55_s_fa1), .B(stage1_c55_s_fa2), .C(stage1_c55_s_fa3), .So(stage2_c55_s_fa5), .Co(stage2_c55_c_fa5));
    FA fa_1246(.A(stage1_c55_s_fa4), .B(stage1_c55_s_fa5), .C(stage1_c55_s_fa6), .So(stage2_c55_s_fa6), .Co(stage2_c55_c_fa6));
    FA fa_1247(.A(stage1_c55_s_fa7), .B(stage1_c55_s_fa8), .C(stage1_c55_s_fa9), .So(stage2_c55_s_fa7), .Co(stage2_c55_c_fa7));
    FA fa_1248(.A(stage1_c55_s_fa10), .B(stage1_c55_s_fa11), .C(stage1_c55_s_fa12), .So(stage2_c55_s_fa8), .Co(stage2_c55_c_fa8));
    FA fa_1249(.A(stage1_c55_c_fa0), .B(stage1_c55_c_fa1), .C(stage1_c55_c_fa2), .So(stage2_c56_s_fa0), .Co(stage2_c56_c_fa0));
    FA fa_1250(.A(stage1_c55_c_fa3), .B(stage1_c55_c_fa4), .C(stage1_c55_c_fa5), .So(stage2_c56_s_fa1), .Co(stage2_c56_c_fa1));
    FA fa_1251(.A(stage1_c55_c_fa6), .B(stage1_c55_c_fa7), .C(stage1_c55_c_fa8), .So(stage2_c56_s_fa2), .Co(stage2_c56_c_fa2));
    FA fa_1252(.A(stage1_c55_c_fa9), .B(stage1_c55_c_fa10), .C(stage1_c55_c_fa11), .So(stage2_c56_s_fa3), .Co(stage2_c56_c_fa3));
    FA fa_1253(.A(stage1_c55_c_fa12), .B(stage1_c55_c_ha0), .C(stage1_c56_s_fa0), .So(stage2_c56_s_fa4), .Co(stage2_c56_c_fa4));
    FA fa_1254(.A(stage1_c56_s_fa1), .B(stage1_c56_s_fa2), .C(stage1_c56_s_fa3), .So(stage2_c56_s_fa5), .Co(stage2_c56_c_fa5));
    FA fa_1255(.A(stage1_c56_s_fa4), .B(stage1_c56_s_fa5), .C(stage1_c56_s_fa6), .So(stage2_c56_s_fa6), .Co(stage2_c56_c_fa6));
    FA fa_1256(.A(stage1_c56_s_fa7), .B(stage1_c56_s_fa8), .C(stage1_c56_s_fa9), .So(stage2_c56_s_fa7), .Co(stage2_c56_c_fa7));
    FA fa_1257(.A(stage1_c56_s_fa10), .B(stage1_c56_s_fa11), .C(stage1_c56_s_fa12), .So(stage2_c56_s_fa8), .Co(stage2_c56_c_fa8));
    FA fa_1258(.A(stage1_c56_c_fa0), .B(stage1_c56_c_fa1), .C(stage1_c56_c_fa2), .So(stage2_c57_s_fa0), .Co(stage2_c57_c_fa0));
    FA fa_1259(.A(stage1_c56_c_fa3), .B(stage1_c56_c_fa4), .C(stage1_c56_c_fa5), .So(stage2_c57_s_fa1), .Co(stage2_c57_c_fa1));
    FA fa_1260(.A(stage1_c56_c_fa6), .B(stage1_c56_c_fa7), .C(stage1_c56_c_fa8), .So(stage2_c57_s_fa2), .Co(stage2_c57_c_fa2));
    FA fa_1261(.A(stage1_c56_c_fa9), .B(stage1_c56_c_fa10), .C(stage1_c56_c_fa11), .So(stage2_c57_s_fa3), .Co(stage2_c57_c_fa3));
    FA fa_1262(.A(stage1_c56_c_fa12), .B(stage1_c56_c_ha0), .C(stage1_c57_s_fa0), .So(stage2_c57_s_fa4), .Co(stage2_c57_c_fa4));
    FA fa_1263(.A(stage1_c57_s_fa1), .B(stage1_c57_s_fa2), .C(stage1_c57_s_fa3), .So(stage2_c57_s_fa5), .Co(stage2_c57_c_fa5));
    FA fa_1264(.A(stage1_c57_s_fa4), .B(stage1_c57_s_fa5), .C(stage1_c57_s_fa6), .So(stage2_c57_s_fa6), .Co(stage2_c57_c_fa6));
    FA fa_1265(.A(stage1_c57_s_fa7), .B(stage1_c57_s_fa8), .C(stage1_c57_s_fa9), .So(stage2_c57_s_fa7), .Co(stage2_c57_c_fa7));
    FA fa_1266(.A(stage1_c57_s_fa10), .B(stage1_c57_s_fa11), .C(stage1_c57_s_fa12), .So(stage2_c57_s_fa8), .Co(stage2_c57_c_fa8));
    FA fa_1267(.A(stage1_c57_c_fa0), .B(stage1_c57_c_fa1), .C(stage1_c57_c_fa2), .So(stage2_c58_s_fa0), .Co(stage2_c58_c_fa0));
    FA fa_1268(.A(stage1_c57_c_fa3), .B(stage1_c57_c_fa4), .C(stage1_c57_c_fa5), .So(stage2_c58_s_fa1), .Co(stage2_c58_c_fa1));
    FA fa_1269(.A(stage1_c57_c_fa6), .B(stage1_c57_c_fa7), .C(stage1_c57_c_fa8), .So(stage2_c58_s_fa2), .Co(stage2_c58_c_fa2));
    FA fa_1270(.A(stage1_c57_c_fa9), .B(stage1_c57_c_fa10), .C(stage1_c57_c_fa11), .So(stage2_c58_s_fa3), .Co(stage2_c58_c_fa3));
    FA fa_1271(.A(stage1_c57_c_fa12), .B(stage1_c57_c_ha0), .C(stage1_c58_s_fa0), .So(stage2_c58_s_fa4), .Co(stage2_c58_c_fa4));
    FA fa_1272(.A(stage1_c58_s_fa1), .B(stage1_c58_s_fa2), .C(stage1_c58_s_fa3), .So(stage2_c58_s_fa5), .Co(stage2_c58_c_fa5));
    FA fa_1273(.A(stage1_c58_s_fa4), .B(stage1_c58_s_fa5), .C(stage1_c58_s_fa6), .So(stage2_c58_s_fa6), .Co(stage2_c58_c_fa6));
    FA fa_1274(.A(stage1_c58_s_fa7), .B(stage1_c58_s_fa8), .C(stage1_c58_s_fa9), .So(stage2_c58_s_fa7), .Co(stage2_c58_c_fa7));
    FA fa_1275(.A(stage1_c58_s_fa10), .B(stage1_c58_s_fa11), .C(stage1_c58_s_fa12), .So(stage2_c58_s_fa8), .Co(stage2_c58_c_fa8));
    FA fa_1276(.A(stage1_c58_c_fa0), .B(stage1_c58_c_fa1), .C(stage1_c58_c_fa2), .So(stage2_c59_s_fa0), .Co(stage2_c59_c_fa0));
    FA fa_1277(.A(stage1_c58_c_fa3), .B(stage1_c58_c_fa4), .C(stage1_c58_c_fa5), .So(stage2_c59_s_fa1), .Co(stage2_c59_c_fa1));
    FA fa_1278(.A(stage1_c58_c_fa6), .B(stage1_c58_c_fa7), .C(stage1_c58_c_fa8), .So(stage2_c59_s_fa2), .Co(stage2_c59_c_fa2));
    FA fa_1279(.A(stage1_c58_c_fa9), .B(stage1_c58_c_fa10), .C(stage1_c58_c_fa11), .So(stage2_c59_s_fa3), .Co(stage2_c59_c_fa3));
    FA fa_1280(.A(stage1_c58_c_fa12), .B(stage1_c58_c_ha0), .C(stage1_c59_s_fa0), .So(stage2_c59_s_fa4), .Co(stage2_c59_c_fa4));
    FA fa_1281(.A(stage1_c59_s_fa1), .B(stage1_c59_s_fa2), .C(stage1_c59_s_fa3), .So(stage2_c59_s_fa5), .Co(stage2_c59_c_fa5));
    FA fa_1282(.A(stage1_c59_s_fa4), .B(stage1_c59_s_fa5), .C(stage1_c59_s_fa6), .So(stage2_c59_s_fa6), .Co(stage2_c59_c_fa6));
    FA fa_1283(.A(stage1_c59_s_fa7), .B(stage1_c59_s_fa8), .C(stage1_c59_s_fa9), .So(stage2_c59_s_fa7), .Co(stage2_c59_c_fa7));
    FA fa_1284(.A(stage1_c59_s_fa10), .B(stage1_c59_s_fa11), .C(stage1_c59_s_fa12), .So(stage2_c59_s_fa8), .Co(stage2_c59_c_fa8));
    FA fa_1285(.A(stage1_c59_c_fa0), .B(stage1_c59_c_fa1), .C(stage1_c59_c_fa2), .So(stage2_c60_s_fa0), .Co(stage2_c60_c_fa0));
    FA fa_1286(.A(stage1_c59_c_fa3), .B(stage1_c59_c_fa4), .C(stage1_c59_c_fa5), .So(stage2_c60_s_fa1), .Co(stage2_c60_c_fa1));
    FA fa_1287(.A(stage1_c59_c_fa6), .B(stage1_c59_c_fa7), .C(stage1_c59_c_fa8), .So(stage2_c60_s_fa2), .Co(stage2_c60_c_fa2));
    FA fa_1288(.A(stage1_c59_c_fa9), .B(stage1_c59_c_fa10), .C(stage1_c59_c_fa11), .So(stage2_c60_s_fa3), .Co(stage2_c60_c_fa3));
    FA fa_1289(.A(stage1_c59_c_fa12), .B(stage1_c59_c_ha0), .C(stage1_c60_s_fa0), .So(stage2_c60_s_fa4), .Co(stage2_c60_c_fa4));
    FA fa_1290(.A(stage1_c60_s_fa1), .B(stage1_c60_s_fa2), .C(stage1_c60_s_fa3), .So(stage2_c60_s_fa5), .Co(stage2_c60_c_fa5));
    FA fa_1291(.A(stage1_c60_s_fa4), .B(stage1_c60_s_fa5), .C(stage1_c60_s_fa6), .So(stage2_c60_s_fa6), .Co(stage2_c60_c_fa6));
    FA fa_1292(.A(stage1_c60_s_fa7), .B(stage1_c60_s_fa8), .C(stage1_c60_s_fa9), .So(stage2_c60_s_fa7), .Co(stage2_c60_c_fa7));
    FA fa_1293(.A(stage1_c60_s_fa10), .B(stage1_c60_s_fa11), .C(stage1_c60_s_fa12), .So(stage2_c60_s_fa8), .Co(stage2_c60_c_fa8));
    FA fa_1294(.A(stage1_c60_c_fa0), .B(stage1_c60_c_fa1), .C(stage1_c60_c_fa2), .So(stage2_c61_s_fa0), .Co(stage2_c61_c_fa0));
    FA fa_1295(.A(stage1_c60_c_fa3), .B(stage1_c60_c_fa4), .C(stage1_c60_c_fa5), .So(stage2_c61_s_fa1), .Co(stage2_c61_c_fa1));
    FA fa_1296(.A(stage1_c60_c_fa6), .B(stage1_c60_c_fa7), .C(stage1_c60_c_fa8), .So(stage2_c61_s_fa2), .Co(stage2_c61_c_fa2));
    FA fa_1297(.A(stage1_c60_c_fa9), .B(stage1_c60_c_fa10), .C(stage1_c60_c_fa11), .So(stage2_c61_s_fa3), .Co(stage2_c61_c_fa3));
    FA fa_1298(.A(stage1_c60_c_fa12), .B(stage1_c60_c_ha0), .C(stage1_c61_s_fa0), .So(stage2_c61_s_fa4), .Co(stage2_c61_c_fa4));
    FA fa_1299(.A(stage1_c61_s_fa1), .B(stage1_c61_s_fa2), .C(stage1_c61_s_fa3), .So(stage2_c61_s_fa5), .Co(stage2_c61_c_fa5));
    FA fa_1300(.A(stage1_c61_s_fa4), .B(stage1_c61_s_fa5), .C(stage1_c61_s_fa6), .So(stage2_c61_s_fa6), .Co(stage2_c61_c_fa6));
    FA fa_1301(.A(stage1_c61_s_fa7), .B(stage1_c61_s_fa8), .C(stage1_c61_s_fa9), .So(stage2_c61_s_fa7), .Co(stage2_c61_c_fa7));
    FA fa_1302(.A(stage1_c61_s_fa10), .B(stage1_c61_s_fa11), .C(stage1_c61_s_fa12), .So(stage2_c61_s_fa8), .Co(stage2_c61_c_fa8));
    FA fa_1303(.A(stage1_c61_c_fa0), .B(stage1_c61_c_fa1), .C(stage1_c61_c_fa2), .So(stage2_c62_s_fa0), .Co(stage2_c62_c_fa0));
    FA fa_1304(.A(stage1_c61_c_fa3), .B(stage1_c61_c_fa4), .C(stage1_c61_c_fa5), .So(stage2_c62_s_fa1), .Co(stage2_c62_c_fa1));
    FA fa_1305(.A(stage1_c61_c_fa6), .B(stage1_c61_c_fa7), .C(stage1_c61_c_fa8), .So(stage2_c62_s_fa2), .Co(stage2_c62_c_fa2));
    FA fa_1306(.A(stage1_c61_c_fa9), .B(stage1_c61_c_fa10), .C(stage1_c61_c_fa11), .So(stage2_c62_s_fa3), .Co(stage2_c62_c_fa3));
    FA fa_1307(.A(stage1_c61_c_fa12), .B(stage1_c61_c_ha0), .C(stage1_c62_s_fa0), .So(stage2_c62_s_fa4), .Co(stage2_c62_c_fa4));
    FA fa_1308(.A(stage1_c62_s_fa1), .B(stage1_c62_s_fa2), .C(stage1_c62_s_fa3), .So(stage2_c62_s_fa5), .Co(stage2_c62_c_fa5));
    FA fa_1309(.A(stage1_c62_s_fa4), .B(stage1_c62_s_fa5), .C(stage1_c62_s_fa6), .So(stage2_c62_s_fa6), .Co(stage2_c62_c_fa6));
    FA fa_1310(.A(stage1_c62_s_fa7), .B(stage1_c62_s_fa8), .C(stage1_c62_s_fa9), .So(stage2_c62_s_fa7), .Co(stage2_c62_c_fa7));
    FA fa_1311(.A(stage1_c62_s_fa10), .B(stage1_c62_s_fa11), .C(stage1_c62_s_fa12), .So(stage2_c62_s_fa8), .Co(stage2_c62_c_fa8));
    FA fa_1312(.A(stage1_c62_c_fa0), .B(stage1_c62_c_fa1), .C(stage1_c62_c_fa2), .So(stage2_c63_s_fa0), .Co(stage2_c63_c_fa0));
    FA fa_1313(.A(stage1_c62_c_fa3), .B(stage1_c62_c_fa4), .C(stage1_c62_c_fa5), .So(stage2_c63_s_fa1), .Co(stage2_c63_c_fa1));
    FA fa_1314(.A(stage1_c62_c_fa6), .B(stage1_c62_c_fa7), .C(stage1_c62_c_fa8), .So(stage2_c63_s_fa2), .Co(stage2_c63_c_fa2));
    FA fa_1315(.A(stage1_c62_c_fa9), .B(stage1_c62_c_fa10), .C(stage1_c62_c_fa11), .So(stage2_c63_s_fa3), .Co(stage2_c63_c_fa3));
    FA fa_1316(.A(stage1_c62_c_fa12), .B(stage1_c62_c_ha0), .C(stage1_c63_s_fa0), .So(stage2_c63_s_fa4), .Co(stage2_c63_c_fa4));
    FA fa_1317(.A(stage1_c63_s_fa1), .B(stage1_c63_s_fa2), .C(stage1_c63_s_fa3), .So(stage2_c63_s_fa5), .Co(stage2_c63_c_fa5));
    FA fa_1318(.A(stage1_c63_s_fa4), .B(stage1_c63_s_fa5), .C(stage1_c63_s_fa6), .So(stage2_c63_s_fa6), .Co(stage2_c63_c_fa6));
    FA fa_1319(.A(stage1_c63_s_fa7), .B(stage1_c63_s_fa8), .C(stage1_c63_s_fa9), .So(stage2_c63_s_fa7), .Co(stage2_c63_c_fa7));
    FA fa_1320(.A(stage1_c63_s_fa10), .B(stage1_c63_s_fa11), .C(stage1_c63_s_fa12), .So(stage2_c63_s_fa8), .Co(stage2_c63_c_fa8));
    FA fa_1321(.A(stage1_c63_c_fa0), .B(stage1_c63_c_fa1), .C(stage1_c63_c_fa2), .So(stage2_c64_s_fa0), .Co(stage2_c64_c_fa0));
    FA fa_1322(.A(stage1_c63_c_fa3), .B(stage1_c63_c_fa4), .C(stage1_c63_c_fa5), .So(stage2_c64_s_fa1), .Co(stage2_c64_c_fa1));
    FA fa_1323(.A(stage1_c63_c_fa6), .B(stage1_c63_c_fa7), .C(stage1_c63_c_fa8), .So(stage2_c64_s_fa2), .Co(stage2_c64_c_fa2));
    FA fa_1324(.A(stage1_c63_c_fa9), .B(stage1_c63_c_fa10), .C(stage1_c63_c_fa11), .So(stage2_c64_s_fa3), .Co(stage2_c64_c_fa3));
    FA fa_1325(.A(stage1_c63_c_fa12), .B(stage1_c63_c_ha0), .C(stage1_c64_s_fa0), .So(stage2_c64_s_fa4), .Co(stage2_c64_c_fa4));
    FA fa_1326(.A(stage1_c64_s_fa1), .B(stage1_c64_s_fa2), .C(stage1_c64_s_fa3), .So(stage2_c64_s_fa5), .Co(stage2_c64_c_fa5));
    FA fa_1327(.A(stage1_c64_s_fa4), .B(stage1_c64_s_fa5), .C(stage1_c64_s_fa6), .So(stage2_c64_s_fa6), .Co(stage2_c64_c_fa6));
    FA fa_1328(.A(stage1_c64_s_fa7), .B(stage1_c64_s_fa8), .C(stage1_c64_s_fa9), .So(stage2_c64_s_fa7), .Co(stage2_c64_c_fa7));
    FA fa_1329(.A(stage1_c64_s_fa10), .B(stage1_c64_s_fa11), .C(stage1_c64_s_fa12), .So(stage2_c64_s_fa8), .Co(stage2_c64_c_fa8));
    FA fa_1330(.A(stage1_c64_c_fa0), .B(stage1_c64_c_fa1), .C(stage1_c64_c_fa2), .So(stage2_c65_s_fa0), .Co(stage2_c65_c_fa0));
    FA fa_1331(.A(stage1_c64_c_fa3), .B(stage1_c64_c_fa4), .C(stage1_c64_c_fa5), .So(stage2_c65_s_fa1), .Co(stage2_c65_c_fa1));
    FA fa_1332(.A(stage1_c64_c_fa6), .B(stage1_c64_c_fa7), .C(stage1_c64_c_fa8), .So(stage2_c65_s_fa2), .Co(stage2_c65_c_fa2));
    FA fa_1333(.A(stage1_c64_c_fa9), .B(stage1_c64_c_fa10), .C(stage1_c64_c_fa11), .So(stage2_c65_s_fa3), .Co(stage2_c65_c_fa3));
    FA fa_1334(.A(stage1_c64_c_fa12), .B(stage1_c64_c_ha0), .C(stage1_c65_s_fa0), .So(stage2_c65_s_fa4), .Co(stage2_c65_c_fa4));
    FA fa_1335(.A(stage1_c65_s_fa1), .B(stage1_c65_s_fa2), .C(stage1_c65_s_fa3), .So(stage2_c65_s_fa5), .Co(stage2_c65_c_fa5));
    FA fa_1336(.A(stage1_c65_s_fa4), .B(stage1_c65_s_fa5), .C(stage1_c65_s_fa6), .So(stage2_c65_s_fa6), .Co(stage2_c65_c_fa6));
    FA fa_1337(.A(stage1_c65_s_fa7), .B(stage1_c65_s_fa8), .C(stage1_c65_s_fa9), .So(stage2_c65_s_fa7), .Co(stage2_c65_c_fa7));
    FA fa_1338(.A(stage1_c65_s_fa10), .B(stage1_c65_s_fa11), .C(stage1_c65_s_fa12), .So(stage2_c65_s_fa8), .Co(stage2_c65_c_fa8));
    FA fa_1339(.A(stage1_c65_c_fa0), .B(stage1_c65_c_fa1), .C(stage1_c65_c_fa2), .So(stage2_c66_s_fa0), .Co(stage2_c66_c_fa0));
    FA fa_1340(.A(stage1_c65_c_fa3), .B(stage1_c65_c_fa4), .C(stage1_c65_c_fa5), .So(stage2_c66_s_fa1), .Co(stage2_c66_c_fa1));
    FA fa_1341(.A(stage1_c65_c_fa6), .B(stage1_c65_c_fa7), .C(stage1_c65_c_fa8), .So(stage2_c66_s_fa2), .Co(stage2_c66_c_fa2));
    FA fa_1342(.A(stage1_c65_c_fa9), .B(stage1_c65_c_fa10), .C(stage1_c65_c_fa11), .So(stage2_c66_s_fa3), .Co(stage2_c66_c_fa3));
    FA fa_1343(.A(stage1_c65_c_fa12), .B(stage1_c65_c_ha0), .C(stage1_c66_s_fa0), .So(stage2_c66_s_fa4), .Co(stage2_c66_c_fa4));
    FA fa_1344(.A(stage1_c66_s_fa1), .B(stage1_c66_s_fa2), .C(stage1_c66_s_fa3), .So(stage2_c66_s_fa5), .Co(stage2_c66_c_fa5));
    FA fa_1345(.A(stage1_c66_s_fa4), .B(stage1_c66_s_fa5), .C(stage1_c66_s_fa6), .So(stage2_c66_s_fa6), .Co(stage2_c66_c_fa6));
    FA fa_1346(.A(stage1_c66_s_fa7), .B(stage1_c66_s_fa8), .C(stage1_c66_s_fa9), .So(stage2_c66_s_fa7), .Co(stage2_c66_c_fa7));
    FA fa_1347(.A(stage1_c66_s_fa10), .B(stage1_c66_s_fa11), .C(stage1_c66_s_fa12), .So(stage2_c66_s_fa8), .Co(stage2_c66_c_fa8));
    FA fa_1348(.A(stage1_c66_c_fa0), .B(stage1_c66_c_fa1), .C(stage1_c66_c_fa2), .So(stage2_c67_s_fa0), .Co(stage2_c67_c_fa0));
    FA fa_1349(.A(stage1_c66_c_fa3), .B(stage1_c66_c_fa4), .C(stage1_c66_c_fa5), .So(stage2_c67_s_fa1), .Co(stage2_c67_c_fa1));
    FA fa_1350(.A(stage1_c66_c_fa6), .B(stage1_c66_c_fa7), .C(stage1_c66_c_fa8), .So(stage2_c67_s_fa2), .Co(stage2_c67_c_fa2));
    FA fa_1351(.A(stage1_c66_c_fa9), .B(stage1_c66_c_fa10), .C(stage1_c66_c_fa11), .So(stage2_c67_s_fa3), .Co(stage2_c67_c_fa3));
    FA fa_1352(.A(stage1_c66_c_fa12), .B(stage1_c66_c_ha0), .C(stage1_c67_s_fa0), .So(stage2_c67_s_fa4), .Co(stage2_c67_c_fa4));
    FA fa_1353(.A(stage1_c67_s_fa1), .B(stage1_c67_s_fa2), .C(stage1_c67_s_fa3), .So(stage2_c67_s_fa5), .Co(stage2_c67_c_fa5));
    FA fa_1354(.A(stage1_c67_s_fa4), .B(stage1_c67_s_fa5), .C(stage1_c67_s_fa6), .So(stage2_c67_s_fa6), .Co(stage2_c67_c_fa6));
    FA fa_1355(.A(stage1_c67_s_fa7), .B(stage1_c67_s_fa8), .C(stage1_c67_s_fa9), .So(stage2_c67_s_fa7), .Co(stage2_c67_c_fa7));
    FA fa_1356(.A(stage1_c67_s_fa10), .B(stage1_c67_s_fa11), .C(stage1_c67_s_fa12), .So(stage2_c67_s_fa8), .Co(stage2_c67_c_fa8));
    FA fa_1357(.A(stage1_c67_c_fa0), .B(stage1_c67_c_fa1), .C(stage1_c67_c_fa2), .So(stage2_c68_s_fa0), .Co(stage2_c68_c_fa0));
    FA fa_1358(.A(stage1_c67_c_fa3), .B(stage1_c67_c_fa4), .C(stage1_c67_c_fa5), .So(stage2_c68_s_fa1), .Co(stage2_c68_c_fa1));
    FA fa_1359(.A(stage1_c67_c_fa6), .B(stage1_c67_c_fa7), .C(stage1_c67_c_fa8), .So(stage2_c68_s_fa2), .Co(stage2_c68_c_fa2));
    FA fa_1360(.A(stage1_c67_c_fa9), .B(stage1_c67_c_fa10), .C(stage1_c67_c_fa11), .So(stage2_c68_s_fa3), .Co(stage2_c68_c_fa3));
    FA fa_1361(.A(stage1_c67_c_fa12), .B(stage1_c67_c_ha0), .C(stage1_c68_s_fa0), .So(stage2_c68_s_fa4), .Co(stage2_c68_c_fa4));
    FA fa_1362(.A(stage1_c68_s_fa1), .B(stage1_c68_s_fa2), .C(stage1_c68_s_fa3), .So(stage2_c68_s_fa5), .Co(stage2_c68_c_fa5));
    FA fa_1363(.A(stage1_c68_s_fa4), .B(stage1_c68_s_fa5), .C(stage1_c68_s_fa6), .So(stage2_c68_s_fa6), .Co(stage2_c68_c_fa6));
    FA fa_1364(.A(stage1_c68_s_fa7), .B(stage1_c68_s_fa8), .C(stage1_c68_s_fa9), .So(stage2_c68_s_fa7), .Co(stage2_c68_c_fa7));
    FA fa_1365(.A(stage1_c68_s_fa10), .B(stage1_c68_s_fa11), .C(stage1_c68_s_fa12), .So(stage2_c68_s_fa8), .Co(stage2_c68_c_fa8));
    FA fa_1366(.A(stage1_c68_c_fa0), .B(stage1_c68_c_fa1), .C(stage1_c68_c_fa2), .So(stage2_c69_s_fa0), .Co(stage2_c69_c_fa0));
    FA fa_1367(.A(stage1_c68_c_fa3), .B(stage1_c68_c_fa4), .C(stage1_c68_c_fa5), .So(stage2_c69_s_fa1), .Co(stage2_c69_c_fa1));
    FA fa_1368(.A(stage1_c68_c_fa6), .B(stage1_c68_c_fa7), .C(stage1_c68_c_fa8), .So(stage2_c69_s_fa2), .Co(stage2_c69_c_fa2));
    FA fa_1369(.A(stage1_c68_c_fa9), .B(stage1_c68_c_fa10), .C(stage1_c68_c_fa11), .So(stage2_c69_s_fa3), .Co(stage2_c69_c_fa3));
    FA fa_1370(.A(stage1_c68_c_fa12), .B(stage1_c68_c_ha0), .C(stage1_c69_s_fa0), .So(stage2_c69_s_fa4), .Co(stage2_c69_c_fa4));
    FA fa_1371(.A(stage1_c69_s_fa1), .B(stage1_c69_s_fa2), .C(stage1_c69_s_fa3), .So(stage2_c69_s_fa5), .Co(stage2_c69_c_fa5));
    FA fa_1372(.A(stage1_c69_s_fa4), .B(stage1_c69_s_fa5), .C(stage1_c69_s_fa6), .So(stage2_c69_s_fa6), .Co(stage2_c69_c_fa6));
    FA fa_1373(.A(stage1_c69_s_fa7), .B(stage1_c69_s_fa8), .C(stage1_c69_s_fa9), .So(stage2_c69_s_fa7), .Co(stage2_c69_c_fa7));
    FA fa_1374(.A(stage1_c69_s_fa10), .B(stage1_c69_s_fa11), .C(stage1_c69_s_fa12), .So(stage2_c69_s_fa8), .Co(stage2_c69_c_fa8));
    FA fa_1375(.A(stage1_c69_c_fa0), .B(stage1_c69_c_fa1), .C(stage1_c69_c_fa2), .So(stage2_c70_s_fa0), .Co(stage2_c70_c_fa0));
    FA fa_1376(.A(stage1_c69_c_fa3), .B(stage1_c69_c_fa4), .C(stage1_c69_c_fa5), .So(stage2_c70_s_fa1), .Co(stage2_c70_c_fa1));
    FA fa_1377(.A(stage1_c69_c_fa6), .B(stage1_c69_c_fa7), .C(stage1_c69_c_fa8), .So(stage2_c70_s_fa2), .Co(stage2_c70_c_fa2));
    FA fa_1378(.A(stage1_c69_c_fa9), .B(stage1_c69_c_fa10), .C(stage1_c69_c_fa11), .So(stage2_c70_s_fa3), .Co(stage2_c70_c_fa3));
    FA fa_1379(.A(stage1_c69_c_fa12), .B(stage1_c69_c_ha0), .C(stage1_c70_s_fa0), .So(stage2_c70_s_fa4), .Co(stage2_c70_c_fa4));
    FA fa_1380(.A(stage1_c70_s_fa1), .B(stage1_c70_s_fa2), .C(stage1_c70_s_fa3), .So(stage2_c70_s_fa5), .Co(stage2_c70_c_fa5));
    FA fa_1381(.A(stage1_c70_s_fa4), .B(stage1_c70_s_fa5), .C(stage1_c70_s_fa6), .So(stage2_c70_s_fa6), .Co(stage2_c70_c_fa6));
    FA fa_1382(.A(stage1_c70_s_fa7), .B(stage1_c70_s_fa8), .C(stage1_c70_s_fa9), .So(stage2_c70_s_fa7), .Co(stage2_c70_c_fa7));
    FA fa_1383(.A(stage1_c70_s_fa10), .B(stage1_c70_s_fa11), .C(stage1_c70_s_fa12), .So(stage2_c70_s_fa8), .Co(stage2_c70_c_fa8));
    FA fa_1384(.A(stage1_c70_c_fa0), .B(stage1_c70_c_fa1), .C(stage1_c70_c_fa2), .So(stage2_c71_s_fa0), .Co(stage2_c71_c_fa0));
    FA fa_1385(.A(stage1_c70_c_fa3), .B(stage1_c70_c_fa4), .C(stage1_c70_c_fa5), .So(stage2_c71_s_fa1), .Co(stage2_c71_c_fa1));
    FA fa_1386(.A(stage1_c70_c_fa6), .B(stage1_c70_c_fa7), .C(stage1_c70_c_fa8), .So(stage2_c71_s_fa2), .Co(stage2_c71_c_fa2));
    FA fa_1387(.A(stage1_c70_c_fa9), .B(stage1_c70_c_fa10), .C(stage1_c70_c_fa11), .So(stage2_c71_s_fa3), .Co(stage2_c71_c_fa3));
    FA fa_1388(.A(stage1_c70_c_fa12), .B(stage1_c70_c_ha0), .C(stage1_c71_s_fa0), .So(stage2_c71_s_fa4), .Co(stage2_c71_c_fa4));
    FA fa_1389(.A(stage1_c71_s_fa1), .B(stage1_c71_s_fa2), .C(stage1_c71_s_fa3), .So(stage2_c71_s_fa5), .Co(stage2_c71_c_fa5));
    FA fa_1390(.A(stage1_c71_s_fa4), .B(stage1_c71_s_fa5), .C(stage1_c71_s_fa6), .So(stage2_c71_s_fa6), .Co(stage2_c71_c_fa6));
    FA fa_1391(.A(stage1_c71_s_fa7), .B(stage1_c71_s_fa8), .C(stage1_c71_s_fa9), .So(stage2_c71_s_fa7), .Co(stage2_c71_c_fa7));
    FA fa_1392(.A(stage1_c71_s_fa10), .B(stage1_c71_s_fa11), .C(stage1_c71_s_fa12), .So(stage2_c71_s_fa8), .Co(stage2_c71_c_fa8));
    FA fa_1393(.A(stage1_c71_c_fa0), .B(stage1_c71_c_fa1), .C(stage1_c71_c_fa2), .So(stage2_c72_s_fa0), .Co(stage2_c72_c_fa0));
    FA fa_1394(.A(stage1_c71_c_fa3), .B(stage1_c71_c_fa4), .C(stage1_c71_c_fa5), .So(stage2_c72_s_fa1), .Co(stage2_c72_c_fa1));
    FA fa_1395(.A(stage1_c71_c_fa6), .B(stage1_c71_c_fa7), .C(stage1_c71_c_fa8), .So(stage2_c72_s_fa2), .Co(stage2_c72_c_fa2));
    FA fa_1396(.A(stage1_c71_c_fa9), .B(stage1_c71_c_fa10), .C(stage1_c71_c_fa11), .So(stage2_c72_s_fa3), .Co(stage2_c72_c_fa3));
    FA fa_1397(.A(stage1_c71_c_fa12), .B(stage1_c71_c_ha0), .C(stage1_c72_s_fa0), .So(stage2_c72_s_fa4), .Co(stage2_c72_c_fa4));
    FA fa_1398(.A(stage1_c72_s_fa1), .B(stage1_c72_s_fa2), .C(stage1_c72_s_fa3), .So(stage2_c72_s_fa5), .Co(stage2_c72_c_fa5));
    FA fa_1399(.A(stage1_c72_s_fa4), .B(stage1_c72_s_fa5), .C(stage1_c72_s_fa6), .So(stage2_c72_s_fa6), .Co(stage2_c72_c_fa6));
    FA fa_1400(.A(stage1_c72_s_fa7), .B(stage1_c72_s_fa8), .C(stage1_c72_s_fa9), .So(stage2_c72_s_fa7), .Co(stage2_c72_c_fa7));
    FA fa_1401(.A(stage1_c72_s_fa10), .B(stage1_c72_s_fa11), .C(stage1_c72_s_fa12), .So(stage2_c72_s_fa8), .Co(stage2_c72_c_fa8));
    FA fa_1402(.A(stage1_c72_c_fa0), .B(stage1_c72_c_fa1), .C(stage1_c72_c_fa2), .So(stage2_c73_s_fa0), .Co(stage2_c73_c_fa0));
    FA fa_1403(.A(stage1_c72_c_fa3), .B(stage1_c72_c_fa4), .C(stage1_c72_c_fa5), .So(stage2_c73_s_fa1), .Co(stage2_c73_c_fa1));
    FA fa_1404(.A(stage1_c72_c_fa6), .B(stage1_c72_c_fa7), .C(stage1_c72_c_fa8), .So(stage2_c73_s_fa2), .Co(stage2_c73_c_fa2));
    FA fa_1405(.A(stage1_c72_c_fa9), .B(stage1_c72_c_fa10), .C(stage1_c72_c_fa11), .So(stage2_c73_s_fa3), .Co(stage2_c73_c_fa3));
    FA fa_1406(.A(stage1_c72_c_fa12), .B(stage1_c73_s_fa0), .C(stage1_c73_s_fa1), .So(stage2_c73_s_fa4), .Co(stage2_c73_c_fa4));
    FA fa_1407(.A(stage1_c73_s_fa2), .B(stage1_c73_s_fa3), .C(stage1_c73_s_fa4), .So(stage2_c73_s_fa5), .Co(stage2_c73_c_fa5));
    FA fa_1408(.A(stage1_c73_s_fa5), .B(stage1_c73_s_fa6), .C(stage1_c73_s_fa7), .So(stage2_c73_s_fa6), .Co(stage2_c73_c_fa6));
    FA fa_1409(.A(stage1_c73_s_fa8), .B(stage1_c73_s_fa9), .C(stage1_c73_s_fa10), .So(stage2_c73_s_fa7), .Co(stage2_c73_c_fa7));
    HA ha_71(.A(stage1_c73_s_fa11), .B(stage1_c73_s_fa12), .So(stage2_c73_s_ha0), .Co(stage2_c73_c_ha0));
    FA fa_1410(.A(stage1_c73_c_fa0), .B(stage1_c73_c_fa1), .C(stage1_c73_c_fa2), .So(stage2_c74_s_fa0), .Co(stage2_c74_c_fa0));
    FA fa_1411(.A(stage1_c73_c_fa3), .B(stage1_c73_c_fa4), .C(stage1_c73_c_fa5), .So(stage2_c74_s_fa1), .Co(stage2_c74_c_fa1));
    FA fa_1412(.A(stage1_c73_c_fa6), .B(stage1_c73_c_fa7), .C(stage1_c73_c_fa8), .So(stage2_c74_s_fa2), .Co(stage2_c74_c_fa2));
    FA fa_1413(.A(stage1_c73_c_fa9), .B(stage1_c73_c_fa10), .C(stage1_c73_c_fa11), .So(stage2_c74_s_fa3), .Co(stage2_c74_c_fa3));
    FA fa_1414(.A(stage1_c73_c_fa12), .B(stage1_c74_s_fa0), .C(stage1_c74_s_fa1), .So(stage2_c74_s_fa4), .Co(stage2_c74_c_fa4));
    FA fa_1415(.A(stage1_c74_s_fa2), .B(stage1_c74_s_fa3), .C(stage1_c74_s_fa4), .So(stage2_c74_s_fa5), .Co(stage2_c74_c_fa5));
    FA fa_1416(.A(stage1_c74_s_fa5), .B(stage1_c74_s_fa6), .C(stage1_c74_s_fa7), .So(stage2_c74_s_fa6), .Co(stage2_c74_c_fa6));
    FA fa_1417(.A(stage1_c74_s_fa8), .B(stage1_c74_s_fa9), .C(stage1_c74_s_fa10), .So(stage2_c74_s_fa7), .Co(stage2_c74_c_fa7));
    HA ha_72(.A(stage1_c74_s_fa11), .B(stage1_c74_s_ha0), .So(stage2_c74_s_ha0), .Co(stage2_c74_c_ha0));
    FA fa_1418(.A(stage1_c74_c_fa0), .B(stage1_c74_c_fa1), .C(stage1_c74_c_fa2), .So(stage2_c75_s_fa0), .Co(stage2_c75_c_fa0));
    FA fa_1419(.A(stage1_c74_c_fa3), .B(stage1_c74_c_fa4), .C(stage1_c74_c_fa5), .So(stage2_c75_s_fa1), .Co(stage2_c75_c_fa1));
    FA fa_1420(.A(stage1_c74_c_fa6), .B(stage1_c74_c_fa7), .C(stage1_c74_c_fa8), .So(stage2_c75_s_fa2), .Co(stage2_c75_c_fa2));
    FA fa_1421(.A(stage1_c74_c_fa9), .B(stage1_c74_c_fa10), .C(stage1_c74_c_fa11), .So(stage2_c75_s_fa3), .Co(stage2_c75_c_fa3));
    FA fa_1422(.A(stage1_c74_c_ha0), .B(stage1_c75_s_fa0), .C(stage1_c75_s_fa1), .So(stage2_c75_s_fa4), .Co(stage2_c75_c_fa4));
    FA fa_1423(.A(stage1_c75_s_fa2), .B(stage1_c75_s_fa3), .C(stage1_c75_s_fa4), .So(stage2_c75_s_fa5), .Co(stage2_c75_c_fa5));
    FA fa_1424(.A(stage1_c75_s_fa5), .B(stage1_c75_s_fa6), .C(stage1_c75_s_fa7), .So(stage2_c75_s_fa6), .Co(stage2_c75_c_fa6));
    FA fa_1425(.A(stage1_c75_s_fa8), .B(stage1_c75_s_fa9), .C(stage1_c75_s_fa10), .So(stage2_c75_s_fa7), .Co(stage2_c75_c_fa7));
    HA ha_73(.A(stage1_c75_s_fa11), .B(stage0_r71_c4), .So(stage2_c75_s_ha0), .Co(stage2_c75_c_ha0));
    FA fa_1426(.A(stage1_c75_c_fa0), .B(stage1_c75_c_fa1), .C(stage1_c75_c_fa2), .So(stage2_c76_s_fa0), .Co(stage2_c76_c_fa0));
    FA fa_1427(.A(stage1_c75_c_fa3), .B(stage1_c75_c_fa4), .C(stage1_c75_c_fa5), .So(stage2_c76_s_fa1), .Co(stage2_c76_c_fa1));
    FA fa_1428(.A(stage1_c75_c_fa6), .B(stage1_c75_c_fa7), .C(stage1_c75_c_fa8), .So(stage2_c76_s_fa2), .Co(stage2_c76_c_fa2));
    FA fa_1429(.A(stage1_c75_c_fa9), .B(stage1_c75_c_fa10), .C(stage1_c75_c_fa11), .So(stage2_c76_s_fa3), .Co(stage2_c76_c_fa3));
    FA fa_1430(.A(stage1_c76_s_fa0), .B(stage1_c76_s_fa1), .C(stage1_c76_s_fa2), .So(stage2_c76_s_fa4), .Co(stage2_c76_c_fa4));
    FA fa_1431(.A(stage1_c76_s_fa3), .B(stage1_c76_s_fa4), .C(stage1_c76_s_fa5), .So(stage2_c76_s_fa5), .Co(stage2_c76_c_fa5));
    FA fa_1432(.A(stage1_c76_s_fa6), .B(stage1_c76_s_fa7), .C(stage1_c76_s_fa8), .So(stage2_c76_s_fa6), .Co(stage2_c76_c_fa6));
    FA fa_1433(.A(stage1_c76_s_fa9), .B(stage1_c76_s_fa10), .C(stage1_c76_s_fa11), .So(stage2_c76_s_fa7), .Co(stage2_c76_c_fa7));
    FA fa_1434(.A(stage1_c76_c_fa0), .B(stage1_c76_c_fa1), .C(stage1_c76_c_fa2), .So(stage2_c77_s_fa0), .Co(stage2_c77_c_fa0));
    FA fa_1435(.A(stage1_c76_c_fa3), .B(stage1_c76_c_fa4), .C(stage1_c76_c_fa5), .So(stage2_c77_s_fa1), .Co(stage2_c77_c_fa1));
    FA fa_1436(.A(stage1_c76_c_fa6), .B(stage1_c76_c_fa7), .C(stage1_c76_c_fa8), .So(stage2_c77_s_fa2), .Co(stage2_c77_c_fa2));
    FA fa_1437(.A(stage1_c76_c_fa9), .B(stage1_c76_c_fa10), .C(stage1_c76_c_fa11), .So(stage2_c77_s_fa3), .Co(stage2_c77_c_fa3));
    FA fa_1438(.A(stage1_c77_s_fa0), .B(stage1_c77_s_fa1), .C(stage1_c77_s_fa2), .So(stage2_c77_s_fa4), .Co(stage2_c77_c_fa4));
    FA fa_1439(.A(stage1_c77_s_fa3), .B(stage1_c77_s_fa4), .C(stage1_c77_s_fa5), .So(stage2_c77_s_fa5), .Co(stage2_c77_c_fa5));
    FA fa_1440(.A(stage1_c77_s_fa6), .B(stage1_c77_s_fa7), .C(stage1_c77_s_fa8), .So(stage2_c77_s_fa6), .Co(stage2_c77_c_fa6));
    FA fa_1441(.A(stage1_c77_s_fa9), .B(stage1_c77_s_fa10), .C(stage1_c77_s_ha0), .So(stage2_c77_s_fa7), .Co(stage2_c77_c_fa7));
    FA fa_1442(.A(stage1_c77_c_fa0), .B(stage1_c77_c_fa1), .C(stage1_c77_c_fa2), .So(stage2_c78_s_fa0), .Co(stage2_c78_c_fa0));
    FA fa_1443(.A(stage1_c77_c_fa3), .B(stage1_c77_c_fa4), .C(stage1_c77_c_fa5), .So(stage2_c78_s_fa1), .Co(stage2_c78_c_fa1));
    FA fa_1444(.A(stage1_c77_c_fa6), .B(stage1_c77_c_fa7), .C(stage1_c77_c_fa8), .So(stage2_c78_s_fa2), .Co(stage2_c78_c_fa2));
    FA fa_1445(.A(stage1_c77_c_fa9), .B(stage1_c77_c_fa10), .C(stage1_c77_c_ha0), .So(stage2_c78_s_fa3), .Co(stage2_c78_c_fa3));
    FA fa_1446(.A(stage1_c78_s_fa0), .B(stage1_c78_s_fa1), .C(stage1_c78_s_fa2), .So(stage2_c78_s_fa4), .Co(stage2_c78_c_fa4));
    FA fa_1447(.A(stage1_c78_s_fa3), .B(stage1_c78_s_fa4), .C(stage1_c78_s_fa5), .So(stage2_c78_s_fa5), .Co(stage2_c78_c_fa5));
    FA fa_1448(.A(stage1_c78_s_fa6), .B(stage1_c78_s_fa7), .C(stage1_c78_s_fa8), .So(stage2_c78_s_fa6), .Co(stage2_c78_c_fa6));
    FA fa_1449(.A(stage1_c78_s_fa9), .B(stage1_c78_s_fa10), .C(stage0_r71_c7), .So(stage2_c78_s_fa7), .Co(stage2_c78_c_fa7));
    FA fa_1450(.A(stage1_c78_c_fa0), .B(stage1_c78_c_fa1), .C(stage1_c78_c_fa2), .So(stage2_c79_s_fa0), .Co(stage2_c79_c_fa0));
    FA fa_1451(.A(stage1_c78_c_fa3), .B(stage1_c78_c_fa4), .C(stage1_c78_c_fa5), .So(stage2_c79_s_fa1), .Co(stage2_c79_c_fa1));
    FA fa_1452(.A(stage1_c78_c_fa6), .B(stage1_c78_c_fa7), .C(stage1_c78_c_fa8), .So(stage2_c79_s_fa2), .Co(stage2_c79_c_fa2));
    FA fa_1453(.A(stage1_c78_c_fa9), .B(stage1_c78_c_fa10), .C(stage1_c79_s_fa0), .So(stage2_c79_s_fa3), .Co(stage2_c79_c_fa3));
    FA fa_1454(.A(stage1_c79_s_fa1), .B(stage1_c79_s_fa2), .C(stage1_c79_s_fa3), .So(stage2_c79_s_fa4), .Co(stage2_c79_c_fa4));
    FA fa_1455(.A(stage1_c79_s_fa4), .B(stage1_c79_s_fa5), .C(stage1_c79_s_fa6), .So(stage2_c79_s_fa5), .Co(stage2_c79_c_fa5));
    FA fa_1456(.A(stage1_c79_s_fa7), .B(stage1_c79_s_fa8), .C(stage1_c79_s_fa9), .So(stage2_c79_s_fa6), .Co(stage2_c79_c_fa6));
    FA fa_1457(.A(stage1_c79_c_fa0), .B(stage1_c79_c_fa1), .C(stage1_c79_c_fa2), .So(stage2_c80_s_fa0), .Co(stage2_c80_c_fa0));
    FA fa_1458(.A(stage1_c79_c_fa3), .B(stage1_c79_c_fa4), .C(stage1_c79_c_fa5), .So(stage2_c80_s_fa1), .Co(stage2_c80_c_fa1));
    FA fa_1459(.A(stage1_c79_c_fa6), .B(stage1_c79_c_fa7), .C(stage1_c79_c_fa8), .So(stage2_c80_s_fa2), .Co(stage2_c80_c_fa2));
    FA fa_1460(.A(stage1_c79_c_fa9), .B(stage1_c79_c_fa10), .C(stage1_c80_s_fa0), .So(stage2_c80_s_fa3), .Co(stage2_c80_c_fa3));
    FA fa_1461(.A(stage1_c80_s_fa1), .B(stage1_c80_s_fa2), .C(stage1_c80_s_fa3), .So(stage2_c80_s_fa4), .Co(stage2_c80_c_fa4));
    FA fa_1462(.A(stage1_c80_s_fa4), .B(stage1_c80_s_fa5), .C(stage1_c80_s_fa6), .So(stage2_c80_s_fa5), .Co(stage2_c80_c_fa5));
    FA fa_1463(.A(stage1_c80_s_fa7), .B(stage1_c80_s_fa8), .C(stage1_c80_s_fa9), .So(stage2_c80_s_fa6), .Co(stage2_c80_c_fa6));
    FA fa_1464(.A(stage1_c80_c_fa0), .B(stage1_c80_c_fa1), .C(stage1_c80_c_fa2), .So(stage2_c81_s_fa0), .Co(stage2_c81_c_fa0));
    FA fa_1465(.A(stage1_c80_c_fa3), .B(stage1_c80_c_fa4), .C(stage1_c80_c_fa5), .So(stage2_c81_s_fa1), .Co(stage2_c81_c_fa1));
    FA fa_1466(.A(stage1_c80_c_fa6), .B(stage1_c80_c_fa7), .C(stage1_c80_c_fa8), .So(stage2_c81_s_fa2), .Co(stage2_c81_c_fa2));
    FA fa_1467(.A(stage1_c80_c_fa9), .B(stage1_c80_c_ha0), .C(stage1_c81_s_fa0), .So(stage2_c81_s_fa3), .Co(stage2_c81_c_fa3));
    FA fa_1468(.A(stage1_c81_s_fa1), .B(stage1_c81_s_fa2), .C(stage1_c81_s_fa3), .So(stage2_c81_s_fa4), .Co(stage2_c81_c_fa4));
    FA fa_1469(.A(stage1_c81_s_fa4), .B(stage1_c81_s_fa5), .C(stage1_c81_s_fa6), .So(stage2_c81_s_fa5), .Co(stage2_c81_c_fa5));
    FA fa_1470(.A(stage1_c81_s_fa7), .B(stage1_c81_s_fa8), .C(stage1_c81_s_fa9), .So(stage2_c81_s_fa6), .Co(stage2_c81_c_fa6));
    FA fa_1471(.A(stage1_c81_c_fa0), .B(stage1_c81_c_fa1), .C(stage1_c81_c_fa2), .So(stage2_c82_s_fa0), .Co(stage2_c82_c_fa0));
    FA fa_1472(.A(stage1_c81_c_fa3), .B(stage1_c81_c_fa4), .C(stage1_c81_c_fa5), .So(stage2_c82_s_fa1), .Co(stage2_c82_c_fa1));
    FA fa_1473(.A(stage1_c81_c_fa6), .B(stage1_c81_c_fa7), .C(stage1_c81_c_fa8), .So(stage2_c82_s_fa2), .Co(stage2_c82_c_fa2));
    FA fa_1474(.A(stage1_c81_c_fa9), .B(stage1_c82_s_fa0), .C(stage1_c82_s_fa1), .So(stage2_c82_s_fa3), .Co(stage2_c82_c_fa3));
    FA fa_1475(.A(stage1_c82_s_fa2), .B(stage1_c82_s_fa3), .C(stage1_c82_s_fa4), .So(stage2_c82_s_fa4), .Co(stage2_c82_c_fa4));
    FA fa_1476(.A(stage1_c82_s_fa5), .B(stage1_c82_s_fa6), .C(stage1_c82_s_fa7), .So(stage2_c82_s_fa5), .Co(stage2_c82_c_fa5));
    HA ha_74(.A(stage1_c82_s_fa8), .B(stage1_c82_s_fa9), .So(stage2_c82_s_ha0), .Co(stage2_c82_c_ha0));
    FA fa_1477(.A(stage1_c82_c_fa0), .B(stage1_c82_c_fa1), .C(stage1_c82_c_fa2), .So(stage2_c83_s_fa0), .Co(stage2_c83_c_fa0));
    FA fa_1478(.A(stage1_c82_c_fa3), .B(stage1_c82_c_fa4), .C(stage1_c82_c_fa5), .So(stage2_c83_s_fa1), .Co(stage2_c83_c_fa1));
    FA fa_1479(.A(stage1_c82_c_fa6), .B(stage1_c82_c_fa7), .C(stage1_c82_c_fa8), .So(stage2_c83_s_fa2), .Co(stage2_c83_c_fa2));
    FA fa_1480(.A(stage1_c82_c_fa9), .B(stage1_c83_s_fa0), .C(stage1_c83_s_fa1), .So(stage2_c83_s_fa3), .Co(stage2_c83_c_fa3));
    FA fa_1481(.A(stage1_c83_s_fa2), .B(stage1_c83_s_fa3), .C(stage1_c83_s_fa4), .So(stage2_c83_s_fa4), .Co(stage2_c83_c_fa4));
    FA fa_1482(.A(stage1_c83_s_fa5), .B(stage1_c83_s_fa6), .C(stage1_c83_s_fa7), .So(stage2_c83_s_fa5), .Co(stage2_c83_c_fa5));
    HA ha_75(.A(stage1_c83_s_fa8), .B(stage1_c83_s_ha0), .So(stage2_c83_s_ha0), .Co(stage2_c83_c_ha0));
    FA fa_1483(.A(stage1_c83_c_fa0), .B(stage1_c83_c_fa1), .C(stage1_c83_c_fa2), .So(stage2_c84_s_fa0), .Co(stage2_c84_c_fa0));
    FA fa_1484(.A(stage1_c83_c_fa3), .B(stage1_c83_c_fa4), .C(stage1_c83_c_fa5), .So(stage2_c84_s_fa1), .Co(stage2_c84_c_fa1));
    FA fa_1485(.A(stage1_c83_c_fa6), .B(stage1_c83_c_fa7), .C(stage1_c83_c_fa8), .So(stage2_c84_s_fa2), .Co(stage2_c84_c_fa2));
    FA fa_1486(.A(stage1_c83_c_ha0), .B(stage1_c84_s_fa0), .C(stage1_c84_s_fa1), .So(stage2_c84_s_fa3), .Co(stage2_c84_c_fa3));
    FA fa_1487(.A(stage1_c84_s_fa2), .B(stage1_c84_s_fa3), .C(stage1_c84_s_fa4), .So(stage2_c84_s_fa4), .Co(stage2_c84_c_fa4));
    FA fa_1488(.A(stage1_c84_s_fa5), .B(stage1_c84_s_fa6), .C(stage1_c84_s_fa7), .So(stage2_c84_s_fa5), .Co(stage2_c84_c_fa5));
    HA ha_76(.A(stage1_c84_s_fa8), .B(stage0_r71_c13), .So(stage2_c84_s_ha0), .Co(stage2_c84_c_ha0));
    FA fa_1489(.A(stage1_c84_c_fa0), .B(stage1_c84_c_fa1), .C(stage1_c84_c_fa2), .So(stage2_c85_s_fa0), .Co(stage2_c85_c_fa0));
    FA fa_1490(.A(stage1_c84_c_fa3), .B(stage1_c84_c_fa4), .C(stage1_c84_c_fa5), .So(stage2_c85_s_fa1), .Co(stage2_c85_c_fa1));
    FA fa_1491(.A(stage1_c84_c_fa6), .B(stage1_c84_c_fa7), .C(stage1_c84_c_fa8), .So(stage2_c85_s_fa2), .Co(stage2_c85_c_fa2));
    FA fa_1492(.A(stage1_c85_s_fa0), .B(stage1_c85_s_fa1), .C(stage1_c85_s_fa2), .So(stage2_c85_s_fa3), .Co(stage2_c85_c_fa3));
    FA fa_1493(.A(stage1_c85_s_fa3), .B(stage1_c85_s_fa4), .C(stage1_c85_s_fa5), .So(stage2_c85_s_fa4), .Co(stage2_c85_c_fa4));
    FA fa_1494(.A(stage1_c85_s_fa6), .B(stage1_c85_s_fa7), .C(stage1_c85_s_fa8), .So(stage2_c85_s_fa5), .Co(stage2_c85_c_fa5));
    FA fa_1495(.A(stage1_c85_c_fa0), .B(stage1_c85_c_fa1), .C(stage1_c85_c_fa2), .So(stage2_c86_s_fa0), .Co(stage2_c86_c_fa0));
    FA fa_1496(.A(stage1_c85_c_fa3), .B(stage1_c85_c_fa4), .C(stage1_c85_c_fa5), .So(stage2_c86_s_fa1), .Co(stage2_c86_c_fa1));
    FA fa_1497(.A(stage1_c85_c_fa6), .B(stage1_c85_c_fa7), .C(stage1_c85_c_fa8), .So(stage2_c86_s_fa2), .Co(stage2_c86_c_fa2));
    FA fa_1498(.A(stage1_c86_s_fa0), .B(stage1_c86_s_fa1), .C(stage1_c86_s_fa2), .So(stage2_c86_s_fa3), .Co(stage2_c86_c_fa3));
    FA fa_1499(.A(stage1_c86_s_fa3), .B(stage1_c86_s_fa4), .C(stage1_c86_s_fa5), .So(stage2_c86_s_fa4), .Co(stage2_c86_c_fa4));
    FA fa_1500(.A(stage1_c86_s_fa6), .B(stage1_c86_s_fa7), .C(stage1_c86_s_ha0), .So(stage2_c86_s_fa5), .Co(stage2_c86_c_fa5));
    FA fa_1501(.A(stage1_c86_c_fa0), .B(stage1_c86_c_fa1), .C(stage1_c86_c_fa2), .So(stage2_c87_s_fa0), .Co(stage2_c87_c_fa0));
    FA fa_1502(.A(stage1_c86_c_fa3), .B(stage1_c86_c_fa4), .C(stage1_c86_c_fa5), .So(stage2_c87_s_fa1), .Co(stage2_c87_c_fa1));
    FA fa_1503(.A(stage1_c86_c_fa6), .B(stage1_c86_c_fa7), .C(stage1_c86_c_ha0), .So(stage2_c87_s_fa2), .Co(stage2_c87_c_fa2));
    FA fa_1504(.A(stage1_c87_s_fa0), .B(stage1_c87_s_fa1), .C(stage1_c87_s_fa2), .So(stage2_c87_s_fa3), .Co(stage2_c87_c_fa3));
    FA fa_1505(.A(stage1_c87_s_fa3), .B(stage1_c87_s_fa4), .C(stage1_c87_s_fa5), .So(stage2_c87_s_fa4), .Co(stage2_c87_c_fa4));
    FA fa_1506(.A(stage1_c87_s_fa6), .B(stage1_c87_s_fa7), .C(stage0_r71_c16), .So(stage2_c87_s_fa5), .Co(stage2_c87_c_fa5));
    FA fa_1507(.A(stage1_c87_c_fa0), .B(stage1_c87_c_fa1), .C(stage1_c87_c_fa2), .So(stage2_c88_s_fa0), .Co(stage2_c88_c_fa0));
    FA fa_1508(.A(stage1_c87_c_fa3), .B(stage1_c87_c_fa4), .C(stage1_c87_c_fa5), .So(stage2_c88_s_fa1), .Co(stage2_c88_c_fa1));
    FA fa_1509(.A(stage1_c87_c_fa6), .B(stage1_c87_c_fa7), .C(stage1_c88_s_fa0), .So(stage2_c88_s_fa2), .Co(stage2_c88_c_fa2));
    FA fa_1510(.A(stage1_c88_s_fa1), .B(stage1_c88_s_fa2), .C(stage1_c88_s_fa3), .So(stage2_c88_s_fa3), .Co(stage2_c88_c_fa3));
    FA fa_1511(.A(stage1_c88_s_fa4), .B(stage1_c88_s_fa5), .C(stage1_c88_s_fa6), .So(stage2_c88_s_fa4), .Co(stage2_c88_c_fa4));
    FA fa_1512(.A(stage1_c88_c_fa0), .B(stage1_c88_c_fa1), .C(stage1_c88_c_fa2), .So(stage2_c89_s_fa0), .Co(stage2_c89_c_fa0));
    FA fa_1513(.A(stage1_c88_c_fa3), .B(stage1_c88_c_fa4), .C(stage1_c88_c_fa5), .So(stage2_c89_s_fa1), .Co(stage2_c89_c_fa1));
    FA fa_1514(.A(stage1_c88_c_fa6), .B(stage1_c88_c_fa7), .C(stage1_c89_s_fa0), .So(stage2_c89_s_fa2), .Co(stage2_c89_c_fa2));
    FA fa_1515(.A(stage1_c89_s_fa1), .B(stage1_c89_s_fa2), .C(stage1_c89_s_fa3), .So(stage2_c89_s_fa3), .Co(stage2_c89_c_fa3));
    FA fa_1516(.A(stage1_c89_s_fa4), .B(stage1_c89_s_fa5), .C(stage1_c89_s_fa6), .So(stage2_c89_s_fa4), .Co(stage2_c89_c_fa4));
    FA fa_1517(.A(stage1_c89_c_fa0), .B(stage1_c89_c_fa1), .C(stage1_c89_c_fa2), .So(stage2_c90_s_fa0), .Co(stage2_c90_c_fa0));
    FA fa_1518(.A(stage1_c89_c_fa3), .B(stage1_c89_c_fa4), .C(stage1_c89_c_fa5), .So(stage2_c90_s_fa1), .Co(stage2_c90_c_fa1));
    FA fa_1519(.A(stage1_c89_c_fa6), .B(stage1_c89_c_ha0), .C(stage1_c90_s_fa0), .So(stage2_c90_s_fa2), .Co(stage2_c90_c_fa2));
    FA fa_1520(.A(stage1_c90_s_fa1), .B(stage1_c90_s_fa2), .C(stage1_c90_s_fa3), .So(stage2_c90_s_fa3), .Co(stage2_c90_c_fa3));
    FA fa_1521(.A(stage1_c90_s_fa4), .B(stage1_c90_s_fa5), .C(stage1_c90_s_fa6), .So(stage2_c90_s_fa4), .Co(stage2_c90_c_fa4));
    FA fa_1522(.A(stage1_c90_c_fa0), .B(stage1_c90_c_fa1), .C(stage1_c90_c_fa2), .So(stage2_c91_s_fa0), .Co(stage2_c91_c_fa0));
    FA fa_1523(.A(stage1_c90_c_fa3), .B(stage1_c90_c_fa4), .C(stage1_c90_c_fa5), .So(stage2_c91_s_fa1), .Co(stage2_c91_c_fa1));
    FA fa_1524(.A(stage1_c90_c_fa6), .B(stage1_c91_s_fa0), .C(stage1_c91_s_fa1), .So(stage2_c91_s_fa2), .Co(stage2_c91_c_fa2));
    FA fa_1525(.A(stage1_c91_s_fa2), .B(stage1_c91_s_fa3), .C(stage1_c91_s_fa4), .So(stage2_c91_s_fa3), .Co(stage2_c91_c_fa3));
    HA ha_77(.A(stage1_c91_s_fa5), .B(stage1_c91_s_fa6), .So(stage2_c91_s_ha0), .Co(stage2_c91_c_ha0));
    FA fa_1526(.A(stage1_c91_c_fa0), .B(stage1_c91_c_fa1), .C(stage1_c91_c_fa2), .So(stage2_c92_s_fa0), .Co(stage2_c92_c_fa0));
    FA fa_1527(.A(stage1_c91_c_fa3), .B(stage1_c91_c_fa4), .C(stage1_c91_c_fa5), .So(stage2_c92_s_fa1), .Co(stage2_c92_c_fa1));
    FA fa_1528(.A(stage1_c91_c_fa6), .B(stage1_c92_s_fa0), .C(stage1_c92_s_fa1), .So(stage2_c92_s_fa2), .Co(stage2_c92_c_fa2));
    FA fa_1529(.A(stage1_c92_s_fa2), .B(stage1_c92_s_fa3), .C(stage1_c92_s_fa4), .So(stage2_c92_s_fa3), .Co(stage2_c92_c_fa3));
    HA ha_78(.A(stage1_c92_s_fa5), .B(stage1_c92_s_ha0), .So(stage2_c92_s_ha0), .Co(stage2_c92_c_ha0));
    FA fa_1530(.A(stage1_c92_c_fa0), .B(stage1_c92_c_fa1), .C(stage1_c92_c_fa2), .So(stage2_c93_s_fa0), .Co(stage2_c93_c_fa0));
    FA fa_1531(.A(stage1_c92_c_fa3), .B(stage1_c92_c_fa4), .C(stage1_c92_c_fa5), .So(stage2_c93_s_fa1), .Co(stage2_c93_c_fa1));
    FA fa_1532(.A(stage1_c92_c_ha0), .B(stage1_c93_s_fa0), .C(stage1_c93_s_fa1), .So(stage2_c93_s_fa2), .Co(stage2_c93_c_fa2));
    FA fa_1533(.A(stage1_c93_s_fa2), .B(stage1_c93_s_fa3), .C(stage1_c93_s_fa4), .So(stage2_c93_s_fa3), .Co(stage2_c93_c_fa3));
    HA ha_79(.A(stage1_c93_s_fa5), .B(stage0_r71_c22), .So(stage2_c93_s_ha0), .Co(stage2_c93_c_ha0));
    FA fa_1534(.A(stage1_c93_c_fa0), .B(stage1_c93_c_fa1), .C(stage1_c93_c_fa2), .So(stage2_c94_s_fa0), .Co(stage2_c94_c_fa0));
    FA fa_1535(.A(stage1_c93_c_fa3), .B(stage1_c93_c_fa4), .C(stage1_c93_c_fa5), .So(stage2_c94_s_fa1), .Co(stage2_c94_c_fa1));
    FA fa_1536(.A(stage1_c94_s_fa0), .B(stage1_c94_s_fa1), .C(stage1_c94_s_fa2), .So(stage2_c94_s_fa2), .Co(stage2_c94_c_fa2));
    FA fa_1537(.A(stage1_c94_s_fa3), .B(stage1_c94_s_fa4), .C(stage1_c94_s_fa5), .So(stage2_c94_s_fa3), .Co(stage2_c94_c_fa3));
    FA fa_1538(.A(stage1_c94_c_fa0), .B(stage1_c94_c_fa1), .C(stage1_c94_c_fa2), .So(stage2_c95_s_fa0), .Co(stage2_c95_c_fa0));
    FA fa_1539(.A(stage1_c94_c_fa3), .B(stage1_c94_c_fa4), .C(stage1_c94_c_fa5), .So(stage2_c95_s_fa1), .Co(stage2_c95_c_fa1));
    FA fa_1540(.A(stage1_c95_s_fa0), .B(stage1_c95_s_fa1), .C(stage1_c95_s_fa2), .So(stage2_c95_s_fa2), .Co(stage2_c95_c_fa2));
    FA fa_1541(.A(stage1_c95_s_fa3), .B(stage1_c95_s_fa4), .C(stage1_c95_s_ha0), .So(stage2_c95_s_fa3), .Co(stage2_c95_c_fa3));
    FA fa_1542(.A(stage1_c95_c_fa0), .B(stage1_c95_c_fa1), .C(stage1_c95_c_fa2), .So(stage2_c96_s_fa0), .Co(stage2_c96_c_fa0));
    FA fa_1543(.A(stage1_c95_c_fa3), .B(stage1_c95_c_fa4), .C(stage1_c95_c_ha0), .So(stage2_c96_s_fa1), .Co(stage2_c96_c_fa1));
    FA fa_1544(.A(stage1_c96_s_fa0), .B(stage1_c96_s_fa1), .C(stage1_c96_s_fa2), .So(stage2_c96_s_fa2), .Co(stage2_c96_c_fa2));
    FA fa_1545(.A(stage1_c96_s_fa3), .B(stage1_c96_s_fa4), .C(stage0_r71_c25), .So(stage2_c96_s_fa3), .Co(stage2_c96_c_fa3));
    FA fa_1546(.A(stage1_c96_c_fa0), .B(stage1_c96_c_fa1), .C(stage1_c96_c_fa2), .So(stage2_c97_s_fa0), .Co(stage2_c97_c_fa0));
    FA fa_1547(.A(stage1_c96_c_fa3), .B(stage1_c96_c_fa4), .C(stage1_c97_s_fa0), .So(stage2_c97_s_fa1), .Co(stage2_c97_c_fa1));
    FA fa_1548(.A(stage1_c97_s_fa1), .B(stage1_c97_s_fa2), .C(stage1_c97_s_fa3), .So(stage2_c97_s_fa2), .Co(stage2_c97_c_fa2));
    FA fa_1549(.A(stage1_c97_c_fa0), .B(stage1_c97_c_fa1), .C(stage1_c97_c_fa2), .So(stage2_c98_s_fa0), .Co(stage2_c98_c_fa0));
    FA fa_1550(.A(stage1_c97_c_fa3), .B(stage1_c97_c_fa4), .C(stage1_c98_s_fa0), .So(stage2_c98_s_fa1), .Co(stage2_c98_c_fa1));
    FA fa_1551(.A(stage1_c98_s_fa1), .B(stage1_c98_s_fa2), .C(stage1_c98_s_fa3), .So(stage2_c98_s_fa2), .Co(stage2_c98_c_fa2));
    FA fa_1552(.A(stage1_c98_c_fa0), .B(stage1_c98_c_fa1), .C(stage1_c98_c_fa2), .So(stage2_c99_s_fa0), .Co(stage2_c99_c_fa0));
    FA fa_1553(.A(stage1_c98_c_fa3), .B(stage1_c98_c_ha0), .C(stage1_c99_s_fa0), .So(stage2_c99_s_fa1), .Co(stage2_c99_c_fa1));
    FA fa_1554(.A(stage1_c99_s_fa1), .B(stage1_c99_s_fa2), .C(stage1_c99_s_fa3), .So(stage2_c99_s_fa2), .Co(stage2_c99_c_fa2));
    FA fa_1555(.A(stage1_c99_c_fa0), .B(stage1_c99_c_fa1), .C(stage1_c99_c_fa2), .So(stage2_c100_s_fa0), .Co(stage2_c100_c_fa0));
    FA fa_1556(.A(stage1_c99_c_fa3), .B(stage1_c100_s_fa0), .C(stage1_c100_s_fa1), .So(stage2_c100_s_fa1), .Co(stage2_c100_c_fa1));
    HA ha_80(.A(stage1_c100_s_fa2), .B(stage1_c100_s_fa3), .So(stage2_c100_s_ha0), .Co(stage2_c100_c_ha0));
    FA fa_1557(.A(stage1_c100_c_fa0), .B(stage1_c100_c_fa1), .C(stage1_c100_c_fa2), .So(stage2_c101_s_fa0), .Co(stage2_c101_c_fa0));
    FA fa_1558(.A(stage1_c100_c_fa3), .B(stage1_c101_s_fa0), .C(stage1_c101_s_fa1), .So(stage2_c101_s_fa1), .Co(stage2_c101_c_fa1));
    HA ha_81(.A(stage1_c101_s_fa2), .B(stage1_c101_s_ha0), .So(stage2_c101_s_ha0), .Co(stage2_c101_c_ha0));
    FA fa_1559(.A(stage1_c101_c_fa0), .B(stage1_c101_c_fa1), .C(stage1_c101_c_fa2), .So(stage2_c102_s_fa0), .Co(stage2_c102_c_fa0));
    FA fa_1560(.A(stage1_c101_c_ha0), .B(stage1_c102_s_fa0), .C(stage1_c102_s_fa1), .So(stage2_c102_s_fa1), .Co(stage2_c102_c_fa1));
    HA ha_82(.A(stage1_c102_s_fa2), .B(stage0_r71_c31), .So(stage2_c102_s_ha0), .Co(stage2_c102_c_ha0));
    FA fa_1561(.A(stage1_c102_c_fa0), .B(stage1_c102_c_fa1), .C(stage1_c102_c_fa2), .So(stage2_c103_s_fa0), .Co(stage2_c103_c_fa0));
    FA fa_1562(.A(stage1_c103_s_fa0), .B(stage1_c103_s_fa1), .C(stage1_c103_s_fa2), .So(stage2_c103_s_fa1), .Co(stage2_c103_c_fa1));
    FA fa_1563(.A(stage1_c103_c_fa0), .B(stage1_c103_c_fa1), .C(stage1_c103_c_fa2), .So(stage2_c104_s_fa0), .Co(stage2_c104_c_fa0));
    FA fa_1564(.A(stage1_c104_s_fa0), .B(stage1_c104_s_fa1), .C(stage1_c104_s_ha0), .So(stage2_c104_s_fa1), .Co(stage2_c104_c_fa1));
    FA fa_1565(.A(stage1_c104_c_fa0), .B(stage1_c104_c_fa1), .C(stage1_c104_c_ha0), .So(stage2_c105_s_fa0), .Co(stage2_c105_c_fa0));
    FA fa_1566(.A(stage1_c105_s_fa0), .B(stage1_c105_s_fa1), .C(stage0_r71_c34), .So(stage2_c105_s_fa1), .Co(stage2_c105_c_fa1));
    FA fa_1567(.A(stage1_c105_c_fa0), .B(stage1_c105_c_fa1), .C(stage1_c106_s_fa0), .So(stage2_c106_s_fa0), .Co(stage2_c106_c_fa0));
    FA fa_1568(.A(stage1_c106_c_fa0), .B(stage1_c106_c_fa1), .C(stage1_c107_s_fa0), .So(stage2_c107_s_fa0), .Co(stage2_c107_c_fa0));
    FA fa_1569(.A(stage1_c107_c_fa0), .B(stage1_c107_c_ha0), .C(stage1_c108_s_fa0), .So(stage2_c108_s_fa0), .Co(stage2_c108_c_fa0));
    HA ha_83(.A(stage1_c108_c_fa0), .B(stage1_c109_s_fa0), .So(stage2_c109_s_ha0), .Co(stage2_c109_c_ha0));
    HA ha_84(.A(stage1_c109_c_fa0), .B(stage1_c110_s_ha0), .So(stage2_c110_s_ha0), .Co(stage2_c110_c_ha0));
    HA ha_85(.A(stage1_c110_c_ha0), .B(stage0_r71_c40), .So(stage2_c111_s_ha0), .Co(stage2_c111_c_ha0));
    HA ha_86(.A(stage2_c2_c_ha0), .B(stage2_c3_s_fa0), .So(stage3_c3_s_ha0), .Co(stage3_c3_c_ha0));
    HA ha_87(.A(stage2_c3_c_fa0), .B(stage2_c4_s_fa0), .So(stage3_c4_s_ha0), .Co(stage3_c4_c_ha0));
    FA fa_1570(.A(stage2_c4_c_fa0), .B(stage2_c5_s_fa0), .C(stage1_c5_s_fa1), .So(stage3_c5_s_fa0), .Co(stage3_c5_c_fa0));
    FA fa_1571(.A(stage2_c5_c_fa0), .B(stage2_c6_s_fa0), .C(stage2_c6_s_ha0), .So(stage3_c6_s_fa0), .Co(stage3_c6_c_fa0));
    FA fa_1572(.A(stage2_c6_c_fa0), .B(stage2_c6_c_ha0), .C(stage2_c7_s_fa0), .So(stage3_c7_s_fa0), .Co(stage3_c7_c_fa0));
    FA fa_1573(.A(stage2_c7_c_fa0), .B(stage2_c7_c_ha0), .C(stage2_c8_s_fa0), .So(stage3_c8_s_fa0), .Co(stage3_c8_c_fa0));
    FA fa_1574(.A(stage2_c8_c_fa0), .B(stage2_c8_c_fa1), .C(stage2_c9_s_fa0), .So(stage3_c9_s_fa0), .Co(stage3_c9_c_fa0));
    HA ha_88(.A(stage2_c9_s_fa1), .B(stage0_r9_c0), .So(stage3_c9_s_ha0), .Co(stage3_c9_c_ha0));
    FA fa_1575(.A(stage2_c9_c_fa0), .B(stage2_c9_c_fa1), .C(stage2_c10_s_fa0), .So(stage3_c10_s_fa0), .Co(stage3_c10_c_fa0));
    HA ha_89(.A(stage2_c10_s_fa1), .B(stage1_c10_s_ha0), .So(stage3_c10_s_ha0), .Co(stage3_c10_c_ha0));
    FA fa_1576(.A(stage2_c10_c_fa0), .B(stage2_c10_c_fa1), .C(stage2_c11_s_fa0), .So(stage3_c11_s_fa0), .Co(stage3_c11_c_fa0));
    HA ha_90(.A(stage2_c11_s_fa1), .B(stage2_c11_s_ha0), .So(stage3_c11_s_ha0), .Co(stage3_c11_c_ha0));
    FA fa_1577(.A(stage2_c11_c_fa0), .B(stage2_c11_c_fa1), .C(stage2_c11_c_ha0), .So(stage3_c12_s_fa0), .Co(stage3_c12_c_fa0));
    FA fa_1578(.A(stage2_c12_s_fa0), .B(stage2_c12_s_fa1), .C(stage2_c12_s_fa2), .So(stage3_c12_s_fa1), .Co(stage3_c12_c_fa1));
    FA fa_1579(.A(stage2_c12_c_fa0), .B(stage2_c12_c_fa1), .C(stage2_c12_c_fa2), .So(stage3_c13_s_fa0), .Co(stage3_c13_c_fa0));
    FA fa_1580(.A(stage2_c13_s_fa0), .B(stage2_c13_s_fa1), .C(stage2_c13_s_fa2), .So(stage3_c13_s_fa1), .Co(stage3_c13_c_fa1));
    FA fa_1581(.A(stage2_c13_c_fa0), .B(stage2_c13_c_fa1), .C(stage2_c13_c_fa2), .So(stage3_c14_s_fa0), .Co(stage3_c14_c_fa0));
    FA fa_1582(.A(stage2_c14_s_fa0), .B(stage2_c14_s_fa1), .C(stage2_c14_s_fa2), .So(stage3_c14_s_fa1), .Co(stage3_c14_c_fa1));
    FA fa_1583(.A(stage2_c14_c_fa0), .B(stage2_c14_c_fa1), .C(stage2_c14_c_fa2), .So(stage3_c15_s_fa0), .Co(stage3_c15_c_fa0));
    FA fa_1584(.A(stage2_c15_s_fa0), .B(stage2_c15_s_fa1), .C(stage2_c15_s_fa2), .So(stage3_c15_s_fa1), .Co(stage3_c15_c_fa1));
    FA fa_1585(.A(stage2_c15_c_fa0), .B(stage2_c15_c_fa1), .C(stage2_c15_c_fa2), .So(stage3_c16_s_fa0), .Co(stage3_c16_c_fa0));
    FA fa_1586(.A(stage2_c15_c_ha0), .B(stage2_c16_s_fa0), .C(stage2_c16_s_fa1), .So(stage3_c16_s_fa1), .Co(stage3_c16_c_fa1));
    HA ha_91(.A(stage2_c16_s_fa2), .B(stage2_c16_s_ha0), .So(stage3_c16_s_ha0), .Co(stage3_c16_c_ha0));
    FA fa_1587(.A(stage2_c16_c_fa0), .B(stage2_c16_c_fa1), .C(stage2_c16_c_fa2), .So(stage3_c17_s_fa0), .Co(stage3_c17_c_fa0));
    FA fa_1588(.A(stage2_c16_c_ha0), .B(stage2_c17_s_fa0), .C(stage2_c17_s_fa1), .So(stage3_c17_s_fa1), .Co(stage3_c17_c_fa1));
    HA ha_92(.A(stage2_c17_s_fa2), .B(stage2_c17_s_fa3), .So(stage3_c17_s_ha0), .Co(stage3_c17_c_ha0));
    FA fa_1589(.A(stage2_c17_c_fa0), .B(stage2_c17_c_fa1), .C(stage2_c17_c_fa2), .So(stage3_c18_s_fa0), .Co(stage3_c18_c_fa0));
    FA fa_1590(.A(stage2_c17_c_fa3), .B(stage2_c18_s_fa0), .C(stage2_c18_s_fa1), .So(stage3_c18_s_fa1), .Co(stage3_c18_c_fa1));
    FA fa_1591(.A(stage2_c18_s_fa2), .B(stage2_c18_s_fa3), .C(stage0_r18_c0), .So(stage3_c18_s_fa2), .Co(stage3_c18_c_fa2));
    FA fa_1592(.A(stage2_c18_c_fa0), .B(stage2_c18_c_fa1), .C(stage2_c18_c_fa2), .So(stage3_c19_s_fa0), .Co(stage3_c19_c_fa0));
    FA fa_1593(.A(stage2_c18_c_fa3), .B(stage2_c19_s_fa0), .C(stage2_c19_s_fa1), .So(stage3_c19_s_fa1), .Co(stage3_c19_c_fa1));
    FA fa_1594(.A(stage2_c19_s_fa2), .B(stage2_c19_s_fa3), .C(stage1_c19_s_ha0), .So(stage3_c19_s_fa2), .Co(stage3_c19_c_fa2));
    FA fa_1595(.A(stage2_c19_c_fa0), .B(stage2_c19_c_fa1), .C(stage2_c19_c_fa2), .So(stage3_c20_s_fa0), .Co(stage3_c20_c_fa0));
    FA fa_1596(.A(stage2_c19_c_fa3), .B(stage2_c20_s_fa0), .C(stage2_c20_s_fa1), .So(stage3_c20_s_fa1), .Co(stage3_c20_c_fa1));
    FA fa_1597(.A(stage2_c20_s_fa2), .B(stage2_c20_s_fa3), .C(stage2_c20_s_ha0), .So(stage3_c20_s_fa2), .Co(stage3_c20_c_fa2));
    FA fa_1598(.A(stage2_c20_c_fa0), .B(stage2_c20_c_fa1), .C(stage2_c20_c_fa2), .So(stage3_c21_s_fa0), .Co(stage3_c21_c_fa0));
    FA fa_1599(.A(stage2_c20_c_fa3), .B(stage2_c20_c_ha0), .C(stage2_c21_s_fa0), .So(stage3_c21_s_fa1), .Co(stage3_c21_c_fa1));
    FA fa_1600(.A(stage2_c21_s_fa1), .B(stage2_c21_s_fa2), .C(stage2_c21_s_fa3), .So(stage3_c21_s_fa2), .Co(stage3_c21_c_fa2));
    FA fa_1601(.A(stage2_c21_c_fa0), .B(stage2_c21_c_fa1), .C(stage2_c21_c_fa2), .So(stage3_c22_s_fa0), .Co(stage3_c22_c_fa0));
    FA fa_1602(.A(stage2_c21_c_fa3), .B(stage2_c21_c_fa4), .C(stage2_c22_s_fa0), .So(stage3_c22_s_fa1), .Co(stage3_c22_c_fa1));
    FA fa_1603(.A(stage2_c22_s_fa1), .B(stage2_c22_s_fa2), .C(stage2_c22_s_fa3), .So(stage3_c22_s_fa2), .Co(stage3_c22_c_fa2));
    FA fa_1604(.A(stage2_c22_c_fa0), .B(stage2_c22_c_fa1), .C(stage2_c22_c_fa2), .So(stage3_c23_s_fa0), .Co(stage3_c23_c_fa0));
    FA fa_1605(.A(stage2_c22_c_fa3), .B(stage2_c22_c_fa4), .C(stage2_c23_s_fa0), .So(stage3_c23_s_fa1), .Co(stage3_c23_c_fa1));
    FA fa_1606(.A(stage2_c23_s_fa1), .B(stage2_c23_s_fa2), .C(stage2_c23_s_fa3), .So(stage3_c23_s_fa2), .Co(stage3_c23_c_fa2));
    HA ha_93(.A(stage2_c23_s_fa4), .B(stage1_c23_s_fa7), .So(stage3_c23_s_ha0), .Co(stage3_c23_c_ha0));
    FA fa_1607(.A(stage2_c23_c_fa0), .B(stage2_c23_c_fa1), .C(stage2_c23_c_fa2), .So(stage3_c24_s_fa0), .Co(stage3_c24_c_fa0));
    FA fa_1608(.A(stage2_c23_c_fa3), .B(stage2_c23_c_fa4), .C(stage2_c24_s_fa0), .So(stage3_c24_s_fa1), .Co(stage3_c24_c_fa1));
    FA fa_1609(.A(stage2_c24_s_fa1), .B(stage2_c24_s_fa2), .C(stage2_c24_s_fa3), .So(stage3_c24_s_fa2), .Co(stage3_c24_c_fa2));
    HA ha_94(.A(stage2_c24_s_fa4), .B(stage2_c24_s_ha0), .So(stage3_c24_s_ha0), .Co(stage3_c24_c_ha0));
    FA fa_1610(.A(stage2_c24_c_fa0), .B(stage2_c24_c_fa1), .C(stage2_c24_c_fa2), .So(stage3_c25_s_fa0), .Co(stage3_c25_c_fa0));
    FA fa_1611(.A(stage2_c24_c_fa3), .B(stage2_c24_c_fa4), .C(stage2_c24_c_ha0), .So(stage3_c25_s_fa1), .Co(stage3_c25_c_fa1));
    FA fa_1612(.A(stage2_c25_s_fa0), .B(stage2_c25_s_fa1), .C(stage2_c25_s_fa2), .So(stage3_c25_s_fa2), .Co(stage3_c25_c_fa2));
    FA fa_1613(.A(stage2_c25_s_fa3), .B(stage2_c25_s_fa4), .C(stage2_c25_s_ha0), .So(stage3_c25_s_fa3), .Co(stage3_c25_c_fa3));
    FA fa_1614(.A(stage2_c25_c_fa0), .B(stage2_c25_c_fa1), .C(stage2_c25_c_fa2), .So(stage3_c26_s_fa0), .Co(stage3_c26_c_fa0));
    FA fa_1615(.A(stage2_c25_c_fa3), .B(stage2_c25_c_fa4), .C(stage2_c25_c_ha0), .So(stage3_c26_s_fa1), .Co(stage3_c26_c_fa1));
    FA fa_1616(.A(stage2_c26_s_fa0), .B(stage2_c26_s_fa1), .C(stage2_c26_s_fa2), .So(stage3_c26_s_fa2), .Co(stage3_c26_c_fa2));
    FA fa_1617(.A(stage2_c26_s_fa3), .B(stage2_c26_s_fa4), .C(stage2_c26_s_fa5), .So(stage3_c26_s_fa3), .Co(stage3_c26_c_fa3));
    FA fa_1618(.A(stage2_c26_c_fa0), .B(stage2_c26_c_fa1), .C(stage2_c26_c_fa2), .So(stage3_c27_s_fa0), .Co(stage3_c27_c_fa0));
    FA fa_1619(.A(stage2_c26_c_fa3), .B(stage2_c26_c_fa4), .C(stage2_c26_c_fa5), .So(stage3_c27_s_fa1), .Co(stage3_c27_c_fa1));
    FA fa_1620(.A(stage2_c27_s_fa0), .B(stage2_c27_s_fa1), .C(stage2_c27_s_fa2), .So(stage3_c27_s_fa2), .Co(stage3_c27_c_fa2));
    FA fa_1621(.A(stage2_c27_s_fa3), .B(stage2_c27_s_fa4), .C(stage2_c27_s_fa5), .So(stage3_c27_s_fa3), .Co(stage3_c27_c_fa3));
    FA fa_1622(.A(stage2_c27_c_fa0), .B(stage2_c27_c_fa1), .C(stage2_c27_c_fa2), .So(stage3_c28_s_fa0), .Co(stage3_c28_c_fa0));
    FA fa_1623(.A(stage2_c27_c_fa3), .B(stage2_c27_c_fa4), .C(stage2_c27_c_fa5), .So(stage3_c28_s_fa1), .Co(stage3_c28_c_fa1));
    FA fa_1624(.A(stage2_c28_s_fa0), .B(stage2_c28_s_fa1), .C(stage2_c28_s_fa2), .So(stage3_c28_s_fa2), .Co(stage3_c28_c_fa2));
    FA fa_1625(.A(stage2_c28_s_fa3), .B(stage2_c28_s_fa4), .C(stage2_c28_s_fa5), .So(stage3_c28_s_fa3), .Co(stage3_c28_c_fa3));
    FA fa_1626(.A(stage2_c28_c_fa0), .B(stage2_c28_c_fa1), .C(stage2_c28_c_fa2), .So(stage3_c29_s_fa0), .Co(stage3_c29_c_fa0));
    FA fa_1627(.A(stage2_c28_c_fa3), .B(stage2_c28_c_fa4), .C(stage2_c28_c_fa5), .So(stage3_c29_s_fa1), .Co(stage3_c29_c_fa1));
    FA fa_1628(.A(stage2_c29_s_fa0), .B(stage2_c29_s_fa1), .C(stage2_c29_s_fa2), .So(stage3_c29_s_fa2), .Co(stage3_c29_c_fa2));
    FA fa_1629(.A(stage2_c29_s_fa3), .B(stage2_c29_s_fa4), .C(stage2_c29_s_fa5), .So(stage3_c29_s_fa3), .Co(stage3_c29_c_fa3));
    FA fa_1630(.A(stage2_c29_c_fa0), .B(stage2_c29_c_fa1), .C(stage2_c29_c_fa2), .So(stage3_c30_s_fa0), .Co(stage3_c30_c_fa0));
    FA fa_1631(.A(stage2_c29_c_fa3), .B(stage2_c29_c_fa4), .C(stage2_c29_c_fa5), .So(stage3_c30_s_fa1), .Co(stage3_c30_c_fa1));
    FA fa_1632(.A(stage2_c29_c_ha0), .B(stage2_c30_s_fa0), .C(stage2_c30_s_fa1), .So(stage3_c30_s_fa2), .Co(stage3_c30_c_fa2));
    FA fa_1633(.A(stage2_c30_s_fa2), .B(stage2_c30_s_fa3), .C(stage2_c30_s_fa4), .So(stage3_c30_s_fa3), .Co(stage3_c30_c_fa3));
    HA ha_95(.A(stage2_c30_s_fa5), .B(stage2_c30_s_fa6), .So(stage3_c30_s_ha0), .Co(stage3_c30_c_ha0));
    FA fa_1634(.A(stage2_c30_c_fa0), .B(stage2_c30_c_fa1), .C(stage2_c30_c_fa2), .So(stage3_c31_s_fa0), .Co(stage3_c31_c_fa0));
    FA fa_1635(.A(stage2_c30_c_fa3), .B(stage2_c30_c_fa4), .C(stage2_c30_c_fa5), .So(stage3_c31_s_fa1), .Co(stage3_c31_c_fa1));
    FA fa_1636(.A(stage2_c30_c_fa6), .B(stage2_c31_s_fa0), .C(stage2_c31_s_fa1), .So(stage3_c31_s_fa2), .Co(stage3_c31_c_fa2));
    FA fa_1637(.A(stage2_c31_s_fa2), .B(stage2_c31_s_fa3), .C(stage2_c31_s_fa4), .So(stage3_c31_s_fa3), .Co(stage3_c31_c_fa3));
    HA ha_96(.A(stage2_c31_s_fa5), .B(stage2_c31_s_fa6), .So(stage3_c31_s_ha0), .Co(stage3_c31_c_ha0));
    FA fa_1638(.A(stage2_c31_c_fa0), .B(stage2_c31_c_fa1), .C(stage2_c31_c_fa2), .So(stage3_c32_s_fa0), .Co(stage3_c32_c_fa0));
    FA fa_1639(.A(stage2_c31_c_fa3), .B(stage2_c31_c_fa4), .C(stage2_c31_c_fa5), .So(stage3_c32_s_fa1), .Co(stage3_c32_c_fa1));
    FA fa_1640(.A(stage2_c31_c_fa6), .B(stage2_c32_s_fa0), .C(stage2_c32_s_fa1), .So(stage3_c32_s_fa2), .Co(stage3_c32_c_fa2));
    FA fa_1641(.A(stage2_c32_s_fa2), .B(stage2_c32_s_fa3), .C(stage2_c32_s_fa4), .So(stage3_c32_s_fa3), .Co(stage3_c32_c_fa3));
    FA fa_1642(.A(stage2_c32_s_fa5), .B(stage2_c32_s_fa6), .C(stage1_c32_s_fa10), .So(stage3_c32_s_fa4), .Co(stage3_c32_c_fa4));
    FA fa_1643(.A(stage2_c32_c_fa0), .B(stage2_c32_c_fa1), .C(stage2_c32_c_fa2), .So(stage3_c33_s_fa0), .Co(stage3_c33_c_fa0));
    FA fa_1644(.A(stage2_c32_c_fa3), .B(stage2_c32_c_fa4), .C(stage2_c32_c_fa5), .So(stage3_c33_s_fa1), .Co(stage3_c33_c_fa1));
    FA fa_1645(.A(stage2_c32_c_fa6), .B(stage2_c33_s_fa0), .C(stage2_c33_s_fa1), .So(stage3_c33_s_fa2), .Co(stage3_c33_c_fa2));
    FA fa_1646(.A(stage2_c33_s_fa2), .B(stage2_c33_s_fa3), .C(stage2_c33_s_fa4), .So(stage3_c33_s_fa3), .Co(stage3_c33_c_fa3));
    FA fa_1647(.A(stage2_c33_s_fa5), .B(stage2_c33_s_fa6), .C(stage2_c33_s_ha0), .So(stage3_c33_s_fa4), .Co(stage3_c33_c_fa4));
    FA fa_1648(.A(stage2_c33_c_fa0), .B(stage2_c33_c_fa1), .C(stage2_c33_c_fa2), .So(stage3_c34_s_fa0), .Co(stage3_c34_c_fa0));
    FA fa_1649(.A(stage2_c33_c_fa3), .B(stage2_c33_c_fa4), .C(stage2_c33_c_fa5), .So(stage3_c34_s_fa1), .Co(stage3_c34_c_fa1));
    FA fa_1650(.A(stage2_c33_c_fa6), .B(stage2_c33_c_ha0), .C(stage2_c34_s_fa0), .So(stage3_c34_s_fa2), .Co(stage3_c34_c_fa2));
    FA fa_1651(.A(stage2_c34_s_fa1), .B(stage2_c34_s_fa2), .C(stage2_c34_s_fa3), .So(stage3_c34_s_fa3), .Co(stage3_c34_c_fa3));
    FA fa_1652(.A(stage2_c34_s_fa4), .B(stage2_c34_s_fa5), .C(stage2_c34_s_fa6), .So(stage3_c34_s_fa4), .Co(stage3_c34_c_fa4));
    FA fa_1653(.A(stage2_c34_c_fa0), .B(stage2_c34_c_fa1), .C(stage2_c34_c_fa2), .So(stage3_c35_s_fa0), .Co(stage3_c35_c_fa0));
    FA fa_1654(.A(stage2_c34_c_fa3), .B(stage2_c34_c_fa4), .C(stage2_c34_c_fa5), .So(stage3_c35_s_fa1), .Co(stage3_c35_c_fa1));
    FA fa_1655(.A(stage2_c34_c_fa6), .B(stage2_c34_c_ha0), .C(stage2_c35_s_fa0), .So(stage3_c35_s_fa2), .Co(stage3_c35_c_fa2));
    FA fa_1656(.A(stage2_c35_s_fa1), .B(stage2_c35_s_fa2), .C(stage2_c35_s_fa3), .So(stage3_c35_s_fa3), .Co(stage3_c35_c_fa3));
    FA fa_1657(.A(stage2_c35_s_fa4), .B(stage2_c35_s_fa5), .C(stage2_c35_s_fa6), .So(stage3_c35_s_fa4), .Co(stage3_c35_c_fa4));
    FA fa_1658(.A(stage2_c35_c_fa0), .B(stage2_c35_c_fa1), .C(stage2_c35_c_fa2), .So(stage3_c36_s_fa0), .Co(stage3_c36_c_fa0));
    FA fa_1659(.A(stage2_c35_c_fa3), .B(stage2_c35_c_fa4), .C(stage2_c35_c_fa5), .So(stage3_c36_s_fa1), .Co(stage3_c36_c_fa1));
    FA fa_1660(.A(stage2_c35_c_fa6), .B(stage2_c35_c_fa7), .C(stage2_c36_s_fa0), .So(stage3_c36_s_fa2), .Co(stage3_c36_c_fa2));
    FA fa_1661(.A(stage2_c36_s_fa1), .B(stage2_c36_s_fa2), .C(stage2_c36_s_fa3), .So(stage3_c36_s_fa3), .Co(stage3_c36_c_fa3));
    FA fa_1662(.A(stage2_c36_s_fa4), .B(stage2_c36_s_fa5), .C(stage2_c36_s_fa6), .So(stage3_c36_s_fa4), .Co(stage3_c36_c_fa4));
    HA ha_97(.A(stage2_c36_s_fa7), .B(stage0_r36_c0), .So(stage3_c36_s_ha0), .Co(stage3_c36_c_ha0));
    FA fa_1663(.A(stage2_c36_c_fa0), .B(stage2_c36_c_fa1), .C(stage2_c36_c_fa2), .So(stage3_c37_s_fa0), .Co(stage3_c37_c_fa0));
    FA fa_1664(.A(stage2_c36_c_fa3), .B(stage2_c36_c_fa4), .C(stage2_c36_c_fa5), .So(stage3_c37_s_fa1), .Co(stage3_c37_c_fa1));
    FA fa_1665(.A(stage2_c36_c_fa6), .B(stage2_c36_c_fa7), .C(stage2_c37_s_fa0), .So(stage3_c37_s_fa2), .Co(stage3_c37_c_fa2));
    FA fa_1666(.A(stage2_c37_s_fa1), .B(stage2_c37_s_fa2), .C(stage2_c37_s_fa3), .So(stage3_c37_s_fa3), .Co(stage3_c37_c_fa3));
    FA fa_1667(.A(stage2_c37_s_fa4), .B(stage2_c37_s_fa5), .C(stage2_c37_s_fa6), .So(stage3_c37_s_fa4), .Co(stage3_c37_c_fa4));
    HA ha_98(.A(stage2_c37_s_fa7), .B(stage1_c37_s_ha0), .So(stage3_c37_s_ha0), .Co(stage3_c37_c_ha0));
    FA fa_1668(.A(stage2_c37_c_fa0), .B(stage2_c37_c_fa1), .C(stage2_c37_c_fa2), .So(stage3_c38_s_fa0), .Co(stage3_c38_c_fa0));
    FA fa_1669(.A(stage2_c37_c_fa3), .B(stage2_c37_c_fa4), .C(stage2_c37_c_fa5), .So(stage3_c38_s_fa1), .Co(stage3_c38_c_fa1));
    FA fa_1670(.A(stage2_c37_c_fa6), .B(stage2_c37_c_fa7), .C(stage2_c38_s_fa0), .So(stage3_c38_s_fa2), .Co(stage3_c38_c_fa2));
    FA fa_1671(.A(stage2_c38_s_fa1), .B(stage2_c38_s_fa2), .C(stage2_c38_s_fa3), .So(stage3_c38_s_fa3), .Co(stage3_c38_c_fa3));
    FA fa_1672(.A(stage2_c38_s_fa4), .B(stage2_c38_s_fa5), .C(stage2_c38_s_fa6), .So(stage3_c38_s_fa4), .Co(stage3_c38_c_fa4));
    HA ha_99(.A(stage2_c38_s_fa7), .B(stage2_c38_s_ha0), .So(stage3_c38_s_ha0), .Co(stage3_c38_c_ha0));
    FA fa_1673(.A(stage2_c38_c_fa0), .B(stage2_c38_c_fa1), .C(stage2_c38_c_fa2), .So(stage3_c39_s_fa0), .Co(stage3_c39_c_fa0));
    FA fa_1674(.A(stage2_c38_c_fa3), .B(stage2_c38_c_fa4), .C(stage2_c38_c_fa5), .So(stage3_c39_s_fa1), .Co(stage3_c39_c_fa1));
    FA fa_1675(.A(stage2_c38_c_fa6), .B(stage2_c38_c_fa7), .C(stage2_c38_c_ha0), .So(stage3_c39_s_fa2), .Co(stage3_c39_c_fa2));
    FA fa_1676(.A(stage2_c39_s_fa0), .B(stage2_c39_s_fa1), .C(stage2_c39_s_fa2), .So(stage3_c39_s_fa3), .Co(stage3_c39_c_fa3));
    FA fa_1677(.A(stage2_c39_s_fa3), .B(stage2_c39_s_fa4), .C(stage2_c39_s_fa5), .So(stage3_c39_s_fa4), .Co(stage3_c39_c_fa4));
    FA fa_1678(.A(stage2_c39_s_fa6), .B(stage2_c39_s_fa7), .C(stage2_c39_s_fa8), .So(stage3_c39_s_fa5), .Co(stage3_c39_c_fa5));
    FA fa_1679(.A(stage2_c39_c_fa0), .B(stage2_c39_c_fa1), .C(stage2_c39_c_fa2), .So(stage3_c40_s_fa0), .Co(stage3_c40_c_fa0));
    FA fa_1680(.A(stage2_c39_c_fa3), .B(stage2_c39_c_fa4), .C(stage2_c39_c_fa5), .So(stage3_c40_s_fa1), .Co(stage3_c40_c_fa1));
    FA fa_1681(.A(stage2_c39_c_fa6), .B(stage2_c39_c_fa7), .C(stage2_c39_c_fa8), .So(stage3_c40_s_fa2), .Co(stage3_c40_c_fa2));
    FA fa_1682(.A(stage2_c40_s_fa0), .B(stage2_c40_s_fa1), .C(stage2_c40_s_fa2), .So(stage3_c40_s_fa3), .Co(stage3_c40_c_fa3));
    FA fa_1683(.A(stage2_c40_s_fa3), .B(stage2_c40_s_fa4), .C(stage2_c40_s_fa5), .So(stage3_c40_s_fa4), .Co(stage3_c40_c_fa4));
    FA fa_1684(.A(stage2_c40_s_fa6), .B(stage2_c40_s_fa7), .C(stage2_c40_s_fa8), .So(stage3_c40_s_fa5), .Co(stage3_c40_c_fa5));
    FA fa_1685(.A(stage2_c40_c_fa0), .B(stage2_c40_c_fa1), .C(stage2_c40_c_fa2), .So(stage3_c41_s_fa0), .Co(stage3_c41_c_fa0));
    FA fa_1686(.A(stage2_c40_c_fa3), .B(stage2_c40_c_fa4), .C(stage2_c40_c_fa5), .So(stage3_c41_s_fa1), .Co(stage3_c41_c_fa1));
    FA fa_1687(.A(stage2_c40_c_fa6), .B(stage2_c40_c_fa7), .C(stage2_c40_c_fa8), .So(stage3_c41_s_fa2), .Co(stage3_c41_c_fa2));
    FA fa_1688(.A(stage2_c41_s_fa0), .B(stage2_c41_s_fa1), .C(stage2_c41_s_fa2), .So(stage3_c41_s_fa3), .Co(stage3_c41_c_fa3));
    FA fa_1689(.A(stage2_c41_s_fa3), .B(stage2_c41_s_fa4), .C(stage2_c41_s_fa5), .So(stage3_c41_s_fa4), .Co(stage3_c41_c_fa4));
    FA fa_1690(.A(stage2_c41_s_fa6), .B(stage2_c41_s_fa7), .C(stage2_c41_s_fa8), .So(stage3_c41_s_fa5), .Co(stage3_c41_c_fa5));
    FA fa_1691(.A(stage2_c41_c_fa0), .B(stage2_c41_c_fa1), .C(stage2_c41_c_fa2), .So(stage3_c42_s_fa0), .Co(stage3_c42_c_fa0));
    FA fa_1692(.A(stage2_c41_c_fa3), .B(stage2_c41_c_fa4), .C(stage2_c41_c_fa5), .So(stage3_c42_s_fa1), .Co(stage3_c42_c_fa1));
    FA fa_1693(.A(stage2_c41_c_fa6), .B(stage2_c41_c_fa7), .C(stage2_c41_c_fa8), .So(stage3_c42_s_fa2), .Co(stage3_c42_c_fa2));
    FA fa_1694(.A(stage2_c42_s_fa0), .B(stage2_c42_s_fa1), .C(stage2_c42_s_fa2), .So(stage3_c42_s_fa3), .Co(stage3_c42_c_fa3));
    FA fa_1695(.A(stage2_c42_s_fa3), .B(stage2_c42_s_fa4), .C(stage2_c42_s_fa5), .So(stage3_c42_s_fa4), .Co(stage3_c42_c_fa4));
    FA fa_1696(.A(stage2_c42_s_fa6), .B(stage2_c42_s_fa7), .C(stage2_c42_s_fa8), .So(stage3_c42_s_fa5), .Co(stage3_c42_c_fa5));
    FA fa_1697(.A(stage2_c42_c_fa0), .B(stage2_c42_c_fa1), .C(stage2_c42_c_fa2), .So(stage3_c43_s_fa0), .Co(stage3_c43_c_fa0));
    FA fa_1698(.A(stage2_c42_c_fa3), .B(stage2_c42_c_fa4), .C(stage2_c42_c_fa5), .So(stage3_c43_s_fa1), .Co(stage3_c43_c_fa1));
    FA fa_1699(.A(stage2_c42_c_fa6), .B(stage2_c42_c_fa7), .C(stage2_c42_c_fa8), .So(stage3_c43_s_fa2), .Co(stage3_c43_c_fa2));
    FA fa_1700(.A(stage2_c43_s_fa0), .B(stage2_c43_s_fa1), .C(stage2_c43_s_fa2), .So(stage3_c43_s_fa3), .Co(stage3_c43_c_fa3));
    FA fa_1701(.A(stage2_c43_s_fa3), .B(stage2_c43_s_fa4), .C(stage2_c43_s_fa5), .So(stage3_c43_s_fa4), .Co(stage3_c43_c_fa4));
    FA fa_1702(.A(stage2_c43_s_fa6), .B(stage2_c43_s_fa7), .C(stage2_c43_s_fa8), .So(stage3_c43_s_fa5), .Co(stage3_c43_c_fa5));
    FA fa_1703(.A(stage2_c43_c_fa0), .B(stage2_c43_c_fa1), .C(stage2_c43_c_fa2), .So(stage3_c44_s_fa0), .Co(stage3_c44_c_fa0));
    FA fa_1704(.A(stage2_c43_c_fa3), .B(stage2_c43_c_fa4), .C(stage2_c43_c_fa5), .So(stage3_c44_s_fa1), .Co(stage3_c44_c_fa1));
    FA fa_1705(.A(stage2_c43_c_fa6), .B(stage2_c43_c_fa7), .C(stage2_c43_c_fa8), .So(stage3_c44_s_fa2), .Co(stage3_c44_c_fa2));
    FA fa_1706(.A(stage2_c44_s_fa0), .B(stage2_c44_s_fa1), .C(stage2_c44_s_fa2), .So(stage3_c44_s_fa3), .Co(stage3_c44_c_fa3));
    FA fa_1707(.A(stage2_c44_s_fa3), .B(stage2_c44_s_fa4), .C(stage2_c44_s_fa5), .So(stage3_c44_s_fa4), .Co(stage3_c44_c_fa4));
    FA fa_1708(.A(stage2_c44_s_fa6), .B(stage2_c44_s_fa7), .C(stage2_c44_s_fa8), .So(stage3_c44_s_fa5), .Co(stage3_c44_c_fa5));
    FA fa_1709(.A(stage2_c44_c_fa0), .B(stage2_c44_c_fa1), .C(stage2_c44_c_fa2), .So(stage3_c45_s_fa0), .Co(stage3_c45_c_fa0));
    FA fa_1710(.A(stage2_c44_c_fa3), .B(stage2_c44_c_fa4), .C(stage2_c44_c_fa5), .So(stage3_c45_s_fa1), .Co(stage3_c45_c_fa1));
    FA fa_1711(.A(stage2_c44_c_fa6), .B(stage2_c44_c_fa7), .C(stage2_c44_c_fa8), .So(stage3_c45_s_fa2), .Co(stage3_c45_c_fa2));
    FA fa_1712(.A(stage2_c45_s_fa0), .B(stage2_c45_s_fa1), .C(stage2_c45_s_fa2), .So(stage3_c45_s_fa3), .Co(stage3_c45_c_fa3));
    FA fa_1713(.A(stage2_c45_s_fa3), .B(stage2_c45_s_fa4), .C(stage2_c45_s_fa5), .So(stage3_c45_s_fa4), .Co(stage3_c45_c_fa4));
    FA fa_1714(.A(stage2_c45_s_fa6), .B(stage2_c45_s_fa7), .C(stage2_c45_s_fa8), .So(stage3_c45_s_fa5), .Co(stage3_c45_c_fa5));
    FA fa_1715(.A(stage2_c45_c_fa0), .B(stage2_c45_c_fa1), .C(stage2_c45_c_fa2), .So(stage3_c46_s_fa0), .Co(stage3_c46_c_fa0));
    FA fa_1716(.A(stage2_c45_c_fa3), .B(stage2_c45_c_fa4), .C(stage2_c45_c_fa5), .So(stage3_c46_s_fa1), .Co(stage3_c46_c_fa1));
    FA fa_1717(.A(stage2_c45_c_fa6), .B(stage2_c45_c_fa7), .C(stage2_c45_c_fa8), .So(stage3_c46_s_fa2), .Co(stage3_c46_c_fa2));
    FA fa_1718(.A(stage2_c46_s_fa0), .B(stage2_c46_s_fa1), .C(stage2_c46_s_fa2), .So(stage3_c46_s_fa3), .Co(stage3_c46_c_fa3));
    FA fa_1719(.A(stage2_c46_s_fa3), .B(stage2_c46_s_fa4), .C(stage2_c46_s_fa5), .So(stage3_c46_s_fa4), .Co(stage3_c46_c_fa4));
    FA fa_1720(.A(stage2_c46_s_fa6), .B(stage2_c46_s_fa7), .C(stage2_c46_s_fa8), .So(stage3_c46_s_fa5), .Co(stage3_c46_c_fa5));
    FA fa_1721(.A(stage2_c46_c_fa0), .B(stage2_c46_c_fa1), .C(stage2_c46_c_fa2), .So(stage3_c47_s_fa0), .Co(stage3_c47_c_fa0));
    FA fa_1722(.A(stage2_c46_c_fa3), .B(stage2_c46_c_fa4), .C(stage2_c46_c_fa5), .So(stage3_c47_s_fa1), .Co(stage3_c47_c_fa1));
    FA fa_1723(.A(stage2_c46_c_fa6), .B(stage2_c46_c_fa7), .C(stage2_c46_c_fa8), .So(stage3_c47_s_fa2), .Co(stage3_c47_c_fa2));
    FA fa_1724(.A(stage2_c47_s_fa0), .B(stage2_c47_s_fa1), .C(stage2_c47_s_fa2), .So(stage3_c47_s_fa3), .Co(stage3_c47_c_fa3));
    FA fa_1725(.A(stage2_c47_s_fa3), .B(stage2_c47_s_fa4), .C(stage2_c47_s_fa5), .So(stage3_c47_s_fa4), .Co(stage3_c47_c_fa4));
    FA fa_1726(.A(stage2_c47_s_fa6), .B(stage2_c47_s_fa7), .C(stage2_c47_s_fa8), .So(stage3_c47_s_fa5), .Co(stage3_c47_c_fa5));
    FA fa_1727(.A(stage2_c47_c_fa0), .B(stage2_c47_c_fa1), .C(stage2_c47_c_fa2), .So(stage3_c48_s_fa0), .Co(stage3_c48_c_fa0));
    FA fa_1728(.A(stage2_c47_c_fa3), .B(stage2_c47_c_fa4), .C(stage2_c47_c_fa5), .So(stage3_c48_s_fa1), .Co(stage3_c48_c_fa1));
    FA fa_1729(.A(stage2_c47_c_fa6), .B(stage2_c47_c_fa7), .C(stage2_c47_c_fa8), .So(stage3_c48_s_fa2), .Co(stage3_c48_c_fa2));
    FA fa_1730(.A(stage2_c48_s_fa0), .B(stage2_c48_s_fa1), .C(stage2_c48_s_fa2), .So(stage3_c48_s_fa3), .Co(stage3_c48_c_fa3));
    FA fa_1731(.A(stage2_c48_s_fa3), .B(stage2_c48_s_fa4), .C(stage2_c48_s_fa5), .So(stage3_c48_s_fa4), .Co(stage3_c48_c_fa4));
    FA fa_1732(.A(stage2_c48_s_fa6), .B(stage2_c48_s_fa7), .C(stage2_c48_s_fa8), .So(stage3_c48_s_fa5), .Co(stage3_c48_c_fa5));
    FA fa_1733(.A(stage2_c48_c_fa0), .B(stage2_c48_c_fa1), .C(stage2_c48_c_fa2), .So(stage3_c49_s_fa0), .Co(stage3_c49_c_fa0));
    FA fa_1734(.A(stage2_c48_c_fa3), .B(stage2_c48_c_fa4), .C(stage2_c48_c_fa5), .So(stage3_c49_s_fa1), .Co(stage3_c49_c_fa1));
    FA fa_1735(.A(stage2_c48_c_fa6), .B(stage2_c48_c_fa7), .C(stage2_c48_c_fa8), .So(stage3_c49_s_fa2), .Co(stage3_c49_c_fa2));
    FA fa_1736(.A(stage2_c49_s_fa0), .B(stage2_c49_s_fa1), .C(stage2_c49_s_fa2), .So(stage3_c49_s_fa3), .Co(stage3_c49_c_fa3));
    FA fa_1737(.A(stage2_c49_s_fa3), .B(stage2_c49_s_fa4), .C(stage2_c49_s_fa5), .So(stage3_c49_s_fa4), .Co(stage3_c49_c_fa4));
    FA fa_1738(.A(stage2_c49_s_fa6), .B(stage2_c49_s_fa7), .C(stage2_c49_s_fa8), .So(stage3_c49_s_fa5), .Co(stage3_c49_c_fa5));
    FA fa_1739(.A(stage2_c49_c_fa0), .B(stage2_c49_c_fa1), .C(stage2_c49_c_fa2), .So(stage3_c50_s_fa0), .Co(stage3_c50_c_fa0));
    FA fa_1740(.A(stage2_c49_c_fa3), .B(stage2_c49_c_fa4), .C(stage2_c49_c_fa5), .So(stage3_c50_s_fa1), .Co(stage3_c50_c_fa1));
    FA fa_1741(.A(stage2_c49_c_fa6), .B(stage2_c49_c_fa7), .C(stage2_c49_c_fa8), .So(stage3_c50_s_fa2), .Co(stage3_c50_c_fa2));
    FA fa_1742(.A(stage2_c50_s_fa0), .B(stage2_c50_s_fa1), .C(stage2_c50_s_fa2), .So(stage3_c50_s_fa3), .Co(stage3_c50_c_fa3));
    FA fa_1743(.A(stage2_c50_s_fa3), .B(stage2_c50_s_fa4), .C(stage2_c50_s_fa5), .So(stage3_c50_s_fa4), .Co(stage3_c50_c_fa4));
    FA fa_1744(.A(stage2_c50_s_fa6), .B(stage2_c50_s_fa7), .C(stage2_c50_s_fa8), .So(stage3_c50_s_fa5), .Co(stage3_c50_c_fa5));
    FA fa_1745(.A(stage2_c50_c_fa0), .B(stage2_c50_c_fa1), .C(stage2_c50_c_fa2), .So(stage3_c51_s_fa0), .Co(stage3_c51_c_fa0));
    FA fa_1746(.A(stage2_c50_c_fa3), .B(stage2_c50_c_fa4), .C(stage2_c50_c_fa5), .So(stage3_c51_s_fa1), .Co(stage3_c51_c_fa1));
    FA fa_1747(.A(stage2_c50_c_fa6), .B(stage2_c50_c_fa7), .C(stage2_c50_c_fa8), .So(stage3_c51_s_fa2), .Co(stage3_c51_c_fa2));
    FA fa_1748(.A(stage2_c51_s_fa0), .B(stage2_c51_s_fa1), .C(stage2_c51_s_fa2), .So(stage3_c51_s_fa3), .Co(stage3_c51_c_fa3));
    FA fa_1749(.A(stage2_c51_s_fa3), .B(stage2_c51_s_fa4), .C(stage2_c51_s_fa5), .So(stage3_c51_s_fa4), .Co(stage3_c51_c_fa4));
    FA fa_1750(.A(stage2_c51_s_fa6), .B(stage2_c51_s_fa7), .C(stage2_c51_s_fa8), .So(stage3_c51_s_fa5), .Co(stage3_c51_c_fa5));
    FA fa_1751(.A(stage2_c51_c_fa0), .B(stage2_c51_c_fa1), .C(stage2_c51_c_fa2), .So(stage3_c52_s_fa0), .Co(stage3_c52_c_fa0));
    FA fa_1752(.A(stage2_c51_c_fa3), .B(stage2_c51_c_fa4), .C(stage2_c51_c_fa5), .So(stage3_c52_s_fa1), .Co(stage3_c52_c_fa1));
    FA fa_1753(.A(stage2_c51_c_fa6), .B(stage2_c51_c_fa7), .C(stage2_c51_c_fa8), .So(stage3_c52_s_fa2), .Co(stage3_c52_c_fa2));
    FA fa_1754(.A(stage2_c52_s_fa0), .B(stage2_c52_s_fa1), .C(stage2_c52_s_fa2), .So(stage3_c52_s_fa3), .Co(stage3_c52_c_fa3));
    FA fa_1755(.A(stage2_c52_s_fa3), .B(stage2_c52_s_fa4), .C(stage2_c52_s_fa5), .So(stage3_c52_s_fa4), .Co(stage3_c52_c_fa4));
    FA fa_1756(.A(stage2_c52_s_fa6), .B(stage2_c52_s_fa7), .C(stage2_c52_s_fa8), .So(stage3_c52_s_fa5), .Co(stage3_c52_c_fa5));
    FA fa_1757(.A(stage2_c52_c_fa0), .B(stage2_c52_c_fa1), .C(stage2_c52_c_fa2), .So(stage3_c53_s_fa0), .Co(stage3_c53_c_fa0));
    FA fa_1758(.A(stage2_c52_c_fa3), .B(stage2_c52_c_fa4), .C(stage2_c52_c_fa5), .So(stage3_c53_s_fa1), .Co(stage3_c53_c_fa1));
    FA fa_1759(.A(stage2_c52_c_fa6), .B(stage2_c52_c_fa7), .C(stage2_c52_c_fa8), .So(stage3_c53_s_fa2), .Co(stage3_c53_c_fa2));
    FA fa_1760(.A(stage2_c53_s_fa0), .B(stage2_c53_s_fa1), .C(stage2_c53_s_fa2), .So(stage3_c53_s_fa3), .Co(stage3_c53_c_fa3));
    FA fa_1761(.A(stage2_c53_s_fa3), .B(stage2_c53_s_fa4), .C(stage2_c53_s_fa5), .So(stage3_c53_s_fa4), .Co(stage3_c53_c_fa4));
    FA fa_1762(.A(stage2_c53_s_fa6), .B(stage2_c53_s_fa7), .C(stage2_c53_s_fa8), .So(stage3_c53_s_fa5), .Co(stage3_c53_c_fa5));
    FA fa_1763(.A(stage2_c53_c_fa0), .B(stage2_c53_c_fa1), .C(stage2_c53_c_fa2), .So(stage3_c54_s_fa0), .Co(stage3_c54_c_fa0));
    FA fa_1764(.A(stage2_c53_c_fa3), .B(stage2_c53_c_fa4), .C(stage2_c53_c_fa5), .So(stage3_c54_s_fa1), .Co(stage3_c54_c_fa1));
    FA fa_1765(.A(stage2_c53_c_fa6), .B(stage2_c53_c_fa7), .C(stage2_c53_c_fa8), .So(stage3_c54_s_fa2), .Co(stage3_c54_c_fa2));
    FA fa_1766(.A(stage2_c54_s_fa0), .B(stage2_c54_s_fa1), .C(stage2_c54_s_fa2), .So(stage3_c54_s_fa3), .Co(stage3_c54_c_fa3));
    FA fa_1767(.A(stage2_c54_s_fa3), .B(stage2_c54_s_fa4), .C(stage2_c54_s_fa5), .So(stage3_c54_s_fa4), .Co(stage3_c54_c_fa4));
    FA fa_1768(.A(stage2_c54_s_fa6), .B(stage2_c54_s_fa7), .C(stage2_c54_s_fa8), .So(stage3_c54_s_fa5), .Co(stage3_c54_c_fa5));
    FA fa_1769(.A(stage2_c54_c_fa0), .B(stage2_c54_c_fa1), .C(stage2_c54_c_fa2), .So(stage3_c55_s_fa0), .Co(stage3_c55_c_fa0));
    FA fa_1770(.A(stage2_c54_c_fa3), .B(stage2_c54_c_fa4), .C(stage2_c54_c_fa5), .So(stage3_c55_s_fa1), .Co(stage3_c55_c_fa1));
    FA fa_1771(.A(stage2_c54_c_fa6), .B(stage2_c54_c_fa7), .C(stage2_c54_c_fa8), .So(stage3_c55_s_fa2), .Co(stage3_c55_c_fa2));
    FA fa_1772(.A(stage2_c55_s_fa0), .B(stage2_c55_s_fa1), .C(stage2_c55_s_fa2), .So(stage3_c55_s_fa3), .Co(stage3_c55_c_fa3));
    FA fa_1773(.A(stage2_c55_s_fa3), .B(stage2_c55_s_fa4), .C(stage2_c55_s_fa5), .So(stage3_c55_s_fa4), .Co(stage3_c55_c_fa4));
    FA fa_1774(.A(stage2_c55_s_fa6), .B(stage2_c55_s_fa7), .C(stage2_c55_s_fa8), .So(stage3_c55_s_fa5), .Co(stage3_c55_c_fa5));
    FA fa_1775(.A(stage2_c55_c_fa0), .B(stage2_c55_c_fa1), .C(stage2_c55_c_fa2), .So(stage3_c56_s_fa0), .Co(stage3_c56_c_fa0));
    FA fa_1776(.A(stage2_c55_c_fa3), .B(stage2_c55_c_fa4), .C(stage2_c55_c_fa5), .So(stage3_c56_s_fa1), .Co(stage3_c56_c_fa1));
    FA fa_1777(.A(stage2_c55_c_fa6), .B(stage2_c55_c_fa7), .C(stage2_c55_c_fa8), .So(stage3_c56_s_fa2), .Co(stage3_c56_c_fa2));
    FA fa_1778(.A(stage2_c56_s_fa0), .B(stage2_c56_s_fa1), .C(stage2_c56_s_fa2), .So(stage3_c56_s_fa3), .Co(stage3_c56_c_fa3));
    FA fa_1779(.A(stage2_c56_s_fa3), .B(stage2_c56_s_fa4), .C(stage2_c56_s_fa5), .So(stage3_c56_s_fa4), .Co(stage3_c56_c_fa4));
    FA fa_1780(.A(stage2_c56_s_fa6), .B(stage2_c56_s_fa7), .C(stage2_c56_s_fa8), .So(stage3_c56_s_fa5), .Co(stage3_c56_c_fa5));
    FA fa_1781(.A(stage2_c56_c_fa0), .B(stage2_c56_c_fa1), .C(stage2_c56_c_fa2), .So(stage3_c57_s_fa0), .Co(stage3_c57_c_fa0));
    FA fa_1782(.A(stage2_c56_c_fa3), .B(stage2_c56_c_fa4), .C(stage2_c56_c_fa5), .So(stage3_c57_s_fa1), .Co(stage3_c57_c_fa1));
    FA fa_1783(.A(stage2_c56_c_fa6), .B(stage2_c56_c_fa7), .C(stage2_c56_c_fa8), .So(stage3_c57_s_fa2), .Co(stage3_c57_c_fa2));
    FA fa_1784(.A(stage2_c57_s_fa0), .B(stage2_c57_s_fa1), .C(stage2_c57_s_fa2), .So(stage3_c57_s_fa3), .Co(stage3_c57_c_fa3));
    FA fa_1785(.A(stage2_c57_s_fa3), .B(stage2_c57_s_fa4), .C(stage2_c57_s_fa5), .So(stage3_c57_s_fa4), .Co(stage3_c57_c_fa4));
    FA fa_1786(.A(stage2_c57_s_fa6), .B(stage2_c57_s_fa7), .C(stage2_c57_s_fa8), .So(stage3_c57_s_fa5), .Co(stage3_c57_c_fa5));
    FA fa_1787(.A(stage2_c57_c_fa0), .B(stage2_c57_c_fa1), .C(stage2_c57_c_fa2), .So(stage3_c58_s_fa0), .Co(stage3_c58_c_fa0));
    FA fa_1788(.A(stage2_c57_c_fa3), .B(stage2_c57_c_fa4), .C(stage2_c57_c_fa5), .So(stage3_c58_s_fa1), .Co(stage3_c58_c_fa1));
    FA fa_1789(.A(stage2_c57_c_fa6), .B(stage2_c57_c_fa7), .C(stage2_c57_c_fa8), .So(stage3_c58_s_fa2), .Co(stage3_c58_c_fa2));
    FA fa_1790(.A(stage2_c58_s_fa0), .B(stage2_c58_s_fa1), .C(stage2_c58_s_fa2), .So(stage3_c58_s_fa3), .Co(stage3_c58_c_fa3));
    FA fa_1791(.A(stage2_c58_s_fa3), .B(stage2_c58_s_fa4), .C(stage2_c58_s_fa5), .So(stage3_c58_s_fa4), .Co(stage3_c58_c_fa4));
    FA fa_1792(.A(stage2_c58_s_fa6), .B(stage2_c58_s_fa7), .C(stage2_c58_s_fa8), .So(stage3_c58_s_fa5), .Co(stage3_c58_c_fa5));
    FA fa_1793(.A(stage2_c58_c_fa0), .B(stage2_c58_c_fa1), .C(stage2_c58_c_fa2), .So(stage3_c59_s_fa0), .Co(stage3_c59_c_fa0));
    FA fa_1794(.A(stage2_c58_c_fa3), .B(stage2_c58_c_fa4), .C(stage2_c58_c_fa5), .So(stage3_c59_s_fa1), .Co(stage3_c59_c_fa1));
    FA fa_1795(.A(stage2_c58_c_fa6), .B(stage2_c58_c_fa7), .C(stage2_c58_c_fa8), .So(stage3_c59_s_fa2), .Co(stage3_c59_c_fa2));
    FA fa_1796(.A(stage2_c59_s_fa0), .B(stage2_c59_s_fa1), .C(stage2_c59_s_fa2), .So(stage3_c59_s_fa3), .Co(stage3_c59_c_fa3));
    FA fa_1797(.A(stage2_c59_s_fa3), .B(stage2_c59_s_fa4), .C(stage2_c59_s_fa5), .So(stage3_c59_s_fa4), .Co(stage3_c59_c_fa4));
    FA fa_1798(.A(stage2_c59_s_fa6), .B(stage2_c59_s_fa7), .C(stage2_c59_s_fa8), .So(stage3_c59_s_fa5), .Co(stage3_c59_c_fa5));
    FA fa_1799(.A(stage2_c59_c_fa0), .B(stage2_c59_c_fa1), .C(stage2_c59_c_fa2), .So(stage3_c60_s_fa0), .Co(stage3_c60_c_fa0));
    FA fa_1800(.A(stage2_c59_c_fa3), .B(stage2_c59_c_fa4), .C(stage2_c59_c_fa5), .So(stage3_c60_s_fa1), .Co(stage3_c60_c_fa1));
    FA fa_1801(.A(stage2_c59_c_fa6), .B(stage2_c59_c_fa7), .C(stage2_c59_c_fa8), .So(stage3_c60_s_fa2), .Co(stage3_c60_c_fa2));
    FA fa_1802(.A(stage2_c60_s_fa0), .B(stage2_c60_s_fa1), .C(stage2_c60_s_fa2), .So(stage3_c60_s_fa3), .Co(stage3_c60_c_fa3));
    FA fa_1803(.A(stage2_c60_s_fa3), .B(stage2_c60_s_fa4), .C(stage2_c60_s_fa5), .So(stage3_c60_s_fa4), .Co(stage3_c60_c_fa4));
    FA fa_1804(.A(stage2_c60_s_fa6), .B(stage2_c60_s_fa7), .C(stage2_c60_s_fa8), .So(stage3_c60_s_fa5), .Co(stage3_c60_c_fa5));
    FA fa_1805(.A(stage2_c60_c_fa0), .B(stage2_c60_c_fa1), .C(stage2_c60_c_fa2), .So(stage3_c61_s_fa0), .Co(stage3_c61_c_fa0));
    FA fa_1806(.A(stage2_c60_c_fa3), .B(stage2_c60_c_fa4), .C(stage2_c60_c_fa5), .So(stage3_c61_s_fa1), .Co(stage3_c61_c_fa1));
    FA fa_1807(.A(stage2_c60_c_fa6), .B(stage2_c60_c_fa7), .C(stage2_c60_c_fa8), .So(stage3_c61_s_fa2), .Co(stage3_c61_c_fa2));
    FA fa_1808(.A(stage2_c61_s_fa0), .B(stage2_c61_s_fa1), .C(stage2_c61_s_fa2), .So(stage3_c61_s_fa3), .Co(stage3_c61_c_fa3));
    FA fa_1809(.A(stage2_c61_s_fa3), .B(stage2_c61_s_fa4), .C(stage2_c61_s_fa5), .So(stage3_c61_s_fa4), .Co(stage3_c61_c_fa4));
    FA fa_1810(.A(stage2_c61_s_fa6), .B(stage2_c61_s_fa7), .C(stage2_c61_s_fa8), .So(stage3_c61_s_fa5), .Co(stage3_c61_c_fa5));
    FA fa_1811(.A(stage2_c61_c_fa0), .B(stage2_c61_c_fa1), .C(stage2_c61_c_fa2), .So(stage3_c62_s_fa0), .Co(stage3_c62_c_fa0));
    FA fa_1812(.A(stage2_c61_c_fa3), .B(stage2_c61_c_fa4), .C(stage2_c61_c_fa5), .So(stage3_c62_s_fa1), .Co(stage3_c62_c_fa1));
    FA fa_1813(.A(stage2_c61_c_fa6), .B(stage2_c61_c_fa7), .C(stage2_c61_c_fa8), .So(stage3_c62_s_fa2), .Co(stage3_c62_c_fa2));
    FA fa_1814(.A(stage2_c62_s_fa0), .B(stage2_c62_s_fa1), .C(stage2_c62_s_fa2), .So(stage3_c62_s_fa3), .Co(stage3_c62_c_fa3));
    FA fa_1815(.A(stage2_c62_s_fa3), .B(stage2_c62_s_fa4), .C(stage2_c62_s_fa5), .So(stage3_c62_s_fa4), .Co(stage3_c62_c_fa4));
    FA fa_1816(.A(stage2_c62_s_fa6), .B(stage2_c62_s_fa7), .C(stage2_c62_s_fa8), .So(stage3_c62_s_fa5), .Co(stage3_c62_c_fa5));
    FA fa_1817(.A(stage2_c62_c_fa0), .B(stage2_c62_c_fa1), .C(stage2_c62_c_fa2), .So(stage3_c63_s_fa0), .Co(stage3_c63_c_fa0));
    FA fa_1818(.A(stage2_c62_c_fa3), .B(stage2_c62_c_fa4), .C(stage2_c62_c_fa5), .So(stage3_c63_s_fa1), .Co(stage3_c63_c_fa1));
    FA fa_1819(.A(stage2_c62_c_fa6), .B(stage2_c62_c_fa7), .C(stage2_c62_c_fa8), .So(stage3_c63_s_fa2), .Co(stage3_c63_c_fa2));
    FA fa_1820(.A(stage2_c63_s_fa0), .B(stage2_c63_s_fa1), .C(stage2_c63_s_fa2), .So(stage3_c63_s_fa3), .Co(stage3_c63_c_fa3));
    FA fa_1821(.A(stage2_c63_s_fa3), .B(stage2_c63_s_fa4), .C(stage2_c63_s_fa5), .So(stage3_c63_s_fa4), .Co(stage3_c63_c_fa4));
    FA fa_1822(.A(stage2_c63_s_fa6), .B(stage2_c63_s_fa7), .C(stage2_c63_s_fa8), .So(stage3_c63_s_fa5), .Co(stage3_c63_c_fa5));
    FA fa_1823(.A(stage2_c63_c_fa0), .B(stage2_c63_c_fa1), .C(stage2_c63_c_fa2), .So(stage3_c64_s_fa0), .Co(stage3_c64_c_fa0));
    FA fa_1824(.A(stage2_c63_c_fa3), .B(stage2_c63_c_fa4), .C(stage2_c63_c_fa5), .So(stage3_c64_s_fa1), .Co(stage3_c64_c_fa1));
    FA fa_1825(.A(stage2_c63_c_fa6), .B(stage2_c63_c_fa7), .C(stage2_c63_c_fa8), .So(stage3_c64_s_fa2), .Co(stage3_c64_c_fa2));
    FA fa_1826(.A(stage2_c64_s_fa0), .B(stage2_c64_s_fa1), .C(stage2_c64_s_fa2), .So(stage3_c64_s_fa3), .Co(stage3_c64_c_fa3));
    FA fa_1827(.A(stage2_c64_s_fa3), .B(stage2_c64_s_fa4), .C(stage2_c64_s_fa5), .So(stage3_c64_s_fa4), .Co(stage3_c64_c_fa4));
    FA fa_1828(.A(stage2_c64_s_fa6), .B(stage2_c64_s_fa7), .C(stage2_c64_s_fa8), .So(stage3_c64_s_fa5), .Co(stage3_c64_c_fa5));
    FA fa_1829(.A(stage2_c64_c_fa0), .B(stage2_c64_c_fa1), .C(stage2_c64_c_fa2), .So(stage3_c65_s_fa0), .Co(stage3_c65_c_fa0));
    FA fa_1830(.A(stage2_c64_c_fa3), .B(stage2_c64_c_fa4), .C(stage2_c64_c_fa5), .So(stage3_c65_s_fa1), .Co(stage3_c65_c_fa1));
    FA fa_1831(.A(stage2_c64_c_fa6), .B(stage2_c64_c_fa7), .C(stage2_c64_c_fa8), .So(stage3_c65_s_fa2), .Co(stage3_c65_c_fa2));
    FA fa_1832(.A(stage2_c65_s_fa0), .B(stage2_c65_s_fa1), .C(stage2_c65_s_fa2), .So(stage3_c65_s_fa3), .Co(stage3_c65_c_fa3));
    FA fa_1833(.A(stage2_c65_s_fa3), .B(stage2_c65_s_fa4), .C(stage2_c65_s_fa5), .So(stage3_c65_s_fa4), .Co(stage3_c65_c_fa4));
    FA fa_1834(.A(stage2_c65_s_fa6), .B(stage2_c65_s_fa7), .C(stage2_c65_s_fa8), .So(stage3_c65_s_fa5), .Co(stage3_c65_c_fa5));
    FA fa_1835(.A(stage2_c65_c_fa0), .B(stage2_c65_c_fa1), .C(stage2_c65_c_fa2), .So(stage3_c66_s_fa0), .Co(stage3_c66_c_fa0));
    FA fa_1836(.A(stage2_c65_c_fa3), .B(stage2_c65_c_fa4), .C(stage2_c65_c_fa5), .So(stage3_c66_s_fa1), .Co(stage3_c66_c_fa1));
    FA fa_1837(.A(stage2_c65_c_fa6), .B(stage2_c65_c_fa7), .C(stage2_c65_c_fa8), .So(stage3_c66_s_fa2), .Co(stage3_c66_c_fa2));
    FA fa_1838(.A(stage2_c66_s_fa0), .B(stage2_c66_s_fa1), .C(stage2_c66_s_fa2), .So(stage3_c66_s_fa3), .Co(stage3_c66_c_fa3));
    FA fa_1839(.A(stage2_c66_s_fa3), .B(stage2_c66_s_fa4), .C(stage2_c66_s_fa5), .So(stage3_c66_s_fa4), .Co(stage3_c66_c_fa4));
    FA fa_1840(.A(stage2_c66_s_fa6), .B(stage2_c66_s_fa7), .C(stage2_c66_s_fa8), .So(stage3_c66_s_fa5), .Co(stage3_c66_c_fa5));
    FA fa_1841(.A(stage2_c66_c_fa0), .B(stage2_c66_c_fa1), .C(stage2_c66_c_fa2), .So(stage3_c67_s_fa0), .Co(stage3_c67_c_fa0));
    FA fa_1842(.A(stage2_c66_c_fa3), .B(stage2_c66_c_fa4), .C(stage2_c66_c_fa5), .So(stage3_c67_s_fa1), .Co(stage3_c67_c_fa1));
    FA fa_1843(.A(stage2_c66_c_fa6), .B(stage2_c66_c_fa7), .C(stage2_c66_c_fa8), .So(stage3_c67_s_fa2), .Co(stage3_c67_c_fa2));
    FA fa_1844(.A(stage2_c67_s_fa0), .B(stage2_c67_s_fa1), .C(stage2_c67_s_fa2), .So(stage3_c67_s_fa3), .Co(stage3_c67_c_fa3));
    FA fa_1845(.A(stage2_c67_s_fa3), .B(stage2_c67_s_fa4), .C(stage2_c67_s_fa5), .So(stage3_c67_s_fa4), .Co(stage3_c67_c_fa4));
    FA fa_1846(.A(stage2_c67_s_fa6), .B(stage2_c67_s_fa7), .C(stage2_c67_s_fa8), .So(stage3_c67_s_fa5), .Co(stage3_c67_c_fa5));
    FA fa_1847(.A(stage2_c67_c_fa0), .B(stage2_c67_c_fa1), .C(stage2_c67_c_fa2), .So(stage3_c68_s_fa0), .Co(stage3_c68_c_fa0));
    FA fa_1848(.A(stage2_c67_c_fa3), .B(stage2_c67_c_fa4), .C(stage2_c67_c_fa5), .So(stage3_c68_s_fa1), .Co(stage3_c68_c_fa1));
    FA fa_1849(.A(stage2_c67_c_fa6), .B(stage2_c67_c_fa7), .C(stage2_c67_c_fa8), .So(stage3_c68_s_fa2), .Co(stage3_c68_c_fa2));
    FA fa_1850(.A(stage2_c68_s_fa0), .B(stage2_c68_s_fa1), .C(stage2_c68_s_fa2), .So(stage3_c68_s_fa3), .Co(stage3_c68_c_fa3));
    FA fa_1851(.A(stage2_c68_s_fa3), .B(stage2_c68_s_fa4), .C(stage2_c68_s_fa5), .So(stage3_c68_s_fa4), .Co(stage3_c68_c_fa4));
    FA fa_1852(.A(stage2_c68_s_fa6), .B(stage2_c68_s_fa7), .C(stage2_c68_s_fa8), .So(stage3_c68_s_fa5), .Co(stage3_c68_c_fa5));
    FA fa_1853(.A(stage2_c68_c_fa0), .B(stage2_c68_c_fa1), .C(stage2_c68_c_fa2), .So(stage3_c69_s_fa0), .Co(stage3_c69_c_fa0));
    FA fa_1854(.A(stage2_c68_c_fa3), .B(stage2_c68_c_fa4), .C(stage2_c68_c_fa5), .So(stage3_c69_s_fa1), .Co(stage3_c69_c_fa1));
    FA fa_1855(.A(stage2_c68_c_fa6), .B(stage2_c68_c_fa7), .C(stage2_c68_c_fa8), .So(stage3_c69_s_fa2), .Co(stage3_c69_c_fa2));
    FA fa_1856(.A(stage2_c69_s_fa0), .B(stage2_c69_s_fa1), .C(stage2_c69_s_fa2), .So(stage3_c69_s_fa3), .Co(stage3_c69_c_fa3));
    FA fa_1857(.A(stage2_c69_s_fa3), .B(stage2_c69_s_fa4), .C(stage2_c69_s_fa5), .So(stage3_c69_s_fa4), .Co(stage3_c69_c_fa4));
    FA fa_1858(.A(stage2_c69_s_fa6), .B(stage2_c69_s_fa7), .C(stage2_c69_s_fa8), .So(stage3_c69_s_fa5), .Co(stage3_c69_c_fa5));
    FA fa_1859(.A(stage2_c69_c_fa0), .B(stage2_c69_c_fa1), .C(stage2_c69_c_fa2), .So(stage3_c70_s_fa0), .Co(stage3_c70_c_fa0));
    FA fa_1860(.A(stage2_c69_c_fa3), .B(stage2_c69_c_fa4), .C(stage2_c69_c_fa5), .So(stage3_c70_s_fa1), .Co(stage3_c70_c_fa1));
    FA fa_1861(.A(stage2_c69_c_fa6), .B(stage2_c69_c_fa7), .C(stage2_c69_c_fa8), .So(stage3_c70_s_fa2), .Co(stage3_c70_c_fa2));
    FA fa_1862(.A(stage2_c70_s_fa0), .B(stage2_c70_s_fa1), .C(stage2_c70_s_fa2), .So(stage3_c70_s_fa3), .Co(stage3_c70_c_fa3));
    FA fa_1863(.A(stage2_c70_s_fa3), .B(stage2_c70_s_fa4), .C(stage2_c70_s_fa5), .So(stage3_c70_s_fa4), .Co(stage3_c70_c_fa4));
    FA fa_1864(.A(stage2_c70_s_fa6), .B(stage2_c70_s_fa7), .C(stage2_c70_s_fa8), .So(stage3_c70_s_fa5), .Co(stage3_c70_c_fa5));
    FA fa_1865(.A(stage2_c70_c_fa0), .B(stage2_c70_c_fa1), .C(stage2_c70_c_fa2), .So(stage3_c71_s_fa0), .Co(stage3_c71_c_fa0));
    FA fa_1866(.A(stage2_c70_c_fa3), .B(stage2_c70_c_fa4), .C(stage2_c70_c_fa5), .So(stage3_c71_s_fa1), .Co(stage3_c71_c_fa1));
    FA fa_1867(.A(stage2_c70_c_fa6), .B(stage2_c70_c_fa7), .C(stage2_c70_c_fa8), .So(stage3_c71_s_fa2), .Co(stage3_c71_c_fa2));
    FA fa_1868(.A(stage2_c71_s_fa0), .B(stage2_c71_s_fa1), .C(stage2_c71_s_fa2), .So(stage3_c71_s_fa3), .Co(stage3_c71_c_fa3));
    FA fa_1869(.A(stage2_c71_s_fa3), .B(stage2_c71_s_fa4), .C(stage2_c71_s_fa5), .So(stage3_c71_s_fa4), .Co(stage3_c71_c_fa4));
    FA fa_1870(.A(stage2_c71_s_fa6), .B(stage2_c71_s_fa7), .C(stage2_c71_s_fa8), .So(stage3_c71_s_fa5), .Co(stage3_c71_c_fa5));
    FA fa_1871(.A(stage2_c71_c_fa0), .B(stage2_c71_c_fa1), .C(stage2_c71_c_fa2), .So(stage3_c72_s_fa0), .Co(stage3_c72_c_fa0));
    FA fa_1872(.A(stage2_c71_c_fa3), .B(stage2_c71_c_fa4), .C(stage2_c71_c_fa5), .So(stage3_c72_s_fa1), .Co(stage3_c72_c_fa1));
    FA fa_1873(.A(stage2_c71_c_fa6), .B(stage2_c71_c_fa7), .C(stage2_c71_c_fa8), .So(stage3_c72_s_fa2), .Co(stage3_c72_c_fa2));
    FA fa_1874(.A(stage2_c72_s_fa0), .B(stage2_c72_s_fa1), .C(stage2_c72_s_fa2), .So(stage3_c72_s_fa3), .Co(stage3_c72_c_fa3));
    FA fa_1875(.A(stage2_c72_s_fa3), .B(stage2_c72_s_fa4), .C(stage2_c72_s_fa5), .So(stage3_c72_s_fa4), .Co(stage3_c72_c_fa4));
    FA fa_1876(.A(stage2_c72_s_fa6), .B(stage2_c72_s_fa7), .C(stage2_c72_s_fa8), .So(stage3_c72_s_fa5), .Co(stage3_c72_c_fa5));
    FA fa_1877(.A(stage2_c72_c_fa0), .B(stage2_c72_c_fa1), .C(stage2_c72_c_fa2), .So(stage3_c73_s_fa0), .Co(stage3_c73_c_fa0));
    FA fa_1878(.A(stage2_c72_c_fa3), .B(stage2_c72_c_fa4), .C(stage2_c72_c_fa5), .So(stage3_c73_s_fa1), .Co(stage3_c73_c_fa1));
    FA fa_1879(.A(stage2_c72_c_fa6), .B(stage2_c72_c_fa7), .C(stage2_c72_c_fa8), .So(stage3_c73_s_fa2), .Co(stage3_c73_c_fa2));
    FA fa_1880(.A(stage2_c73_s_fa0), .B(stage2_c73_s_fa1), .C(stage2_c73_s_fa2), .So(stage3_c73_s_fa3), .Co(stage3_c73_c_fa3));
    FA fa_1881(.A(stage2_c73_s_fa3), .B(stage2_c73_s_fa4), .C(stage2_c73_s_fa5), .So(stage3_c73_s_fa4), .Co(stage3_c73_c_fa4));
    FA fa_1882(.A(stage2_c73_s_fa6), .B(stage2_c73_s_fa7), .C(stage2_c73_s_ha0), .So(stage3_c73_s_fa5), .Co(stage3_c73_c_fa5));
    FA fa_1883(.A(stage2_c73_c_fa0), .B(stage2_c73_c_fa1), .C(stage2_c73_c_fa2), .So(stage3_c74_s_fa0), .Co(stage3_c74_c_fa0));
    FA fa_1884(.A(stage2_c73_c_fa3), .B(stage2_c73_c_fa4), .C(stage2_c73_c_fa5), .So(stage3_c74_s_fa1), .Co(stage3_c74_c_fa1));
    FA fa_1885(.A(stage2_c73_c_fa6), .B(stage2_c73_c_fa7), .C(stage2_c73_c_ha0), .So(stage3_c74_s_fa2), .Co(stage3_c74_c_fa2));
    FA fa_1886(.A(stage2_c74_s_fa0), .B(stage2_c74_s_fa1), .C(stage2_c74_s_fa2), .So(stage3_c74_s_fa3), .Co(stage3_c74_c_fa3));
    FA fa_1887(.A(stage2_c74_s_fa3), .B(stage2_c74_s_fa4), .C(stage2_c74_s_fa5), .So(stage3_c74_s_fa4), .Co(stage3_c74_c_fa4));
    FA fa_1888(.A(stage2_c74_s_fa6), .B(stage2_c74_s_fa7), .C(stage2_c74_s_ha0), .So(stage3_c74_s_fa5), .Co(stage3_c74_c_fa5));
    FA fa_1889(.A(stage2_c74_c_fa0), .B(stage2_c74_c_fa1), .C(stage2_c74_c_fa2), .So(stage3_c75_s_fa0), .Co(stage3_c75_c_fa0));
    FA fa_1890(.A(stage2_c74_c_fa3), .B(stage2_c74_c_fa4), .C(stage2_c74_c_fa5), .So(stage3_c75_s_fa1), .Co(stage3_c75_c_fa1));
    FA fa_1891(.A(stage2_c74_c_fa6), .B(stage2_c74_c_fa7), .C(stage2_c74_c_ha0), .So(stage3_c75_s_fa2), .Co(stage3_c75_c_fa2));
    FA fa_1892(.A(stage2_c75_s_fa0), .B(stage2_c75_s_fa1), .C(stage2_c75_s_fa2), .So(stage3_c75_s_fa3), .Co(stage3_c75_c_fa3));
    FA fa_1893(.A(stage2_c75_s_fa3), .B(stage2_c75_s_fa4), .C(stage2_c75_s_fa5), .So(stage3_c75_s_fa4), .Co(stage3_c75_c_fa4));
    FA fa_1894(.A(stage2_c75_s_fa6), .B(stage2_c75_s_fa7), .C(stage2_c75_s_ha0), .So(stage3_c75_s_fa5), .Co(stage3_c75_c_fa5));
    FA fa_1895(.A(stage2_c75_c_fa0), .B(stage2_c75_c_fa1), .C(stage2_c75_c_fa2), .So(stage3_c76_s_fa0), .Co(stage3_c76_c_fa0));
    FA fa_1896(.A(stage2_c75_c_fa3), .B(stage2_c75_c_fa4), .C(stage2_c75_c_fa5), .So(stage3_c76_s_fa1), .Co(stage3_c76_c_fa1));
    FA fa_1897(.A(stage2_c75_c_fa6), .B(stage2_c75_c_fa7), .C(stage2_c75_c_ha0), .So(stage3_c76_s_fa2), .Co(stage3_c76_c_fa2));
    FA fa_1898(.A(stage2_c76_s_fa0), .B(stage2_c76_s_fa1), .C(stage2_c76_s_fa2), .So(stage3_c76_s_fa3), .Co(stage3_c76_c_fa3));
    FA fa_1899(.A(stage2_c76_s_fa3), .B(stage2_c76_s_fa4), .C(stage2_c76_s_fa5), .So(stage3_c76_s_fa4), .Co(stage3_c76_c_fa4));
    HA ha_100(.A(stage2_c76_s_fa6), .B(stage2_c76_s_fa7), .So(stage3_c76_s_ha0), .Co(stage3_c76_c_ha0));
    FA fa_1900(.A(stage2_c76_c_fa0), .B(stage2_c76_c_fa1), .C(stage2_c76_c_fa2), .So(stage3_c77_s_fa0), .Co(stage3_c77_c_fa0));
    FA fa_1901(.A(stage2_c76_c_fa3), .B(stage2_c76_c_fa4), .C(stage2_c76_c_fa5), .So(stage3_c77_s_fa1), .Co(stage3_c77_c_fa1));
    FA fa_1902(.A(stage2_c76_c_fa6), .B(stage2_c76_c_fa7), .C(stage2_c77_s_fa0), .So(stage3_c77_s_fa2), .Co(stage3_c77_c_fa2));
    FA fa_1903(.A(stage2_c77_s_fa1), .B(stage2_c77_s_fa2), .C(stage2_c77_s_fa3), .So(stage3_c77_s_fa3), .Co(stage3_c77_c_fa3));
    FA fa_1904(.A(stage2_c77_s_fa4), .B(stage2_c77_s_fa5), .C(stage2_c77_s_fa6), .So(stage3_c77_s_fa4), .Co(stage3_c77_c_fa4));
    FA fa_1905(.A(stage2_c77_c_fa0), .B(stage2_c77_c_fa1), .C(stage2_c77_c_fa2), .So(stage3_c78_s_fa0), .Co(stage3_c78_c_fa0));
    FA fa_1906(.A(stage2_c77_c_fa3), .B(stage2_c77_c_fa4), .C(stage2_c77_c_fa5), .So(stage3_c78_s_fa1), .Co(stage3_c78_c_fa1));
    FA fa_1907(.A(stage2_c77_c_fa6), .B(stage2_c77_c_fa7), .C(stage2_c78_s_fa0), .So(stage3_c78_s_fa2), .Co(stage3_c78_c_fa2));
    FA fa_1908(.A(stage2_c78_s_fa1), .B(stage2_c78_s_fa2), .C(stage2_c78_s_fa3), .So(stage3_c78_s_fa3), .Co(stage3_c78_c_fa3));
    FA fa_1909(.A(stage2_c78_s_fa4), .B(stage2_c78_s_fa5), .C(stage2_c78_s_fa6), .So(stage3_c78_s_fa4), .Co(stage3_c78_c_fa4));
    FA fa_1910(.A(stage2_c78_c_fa0), .B(stage2_c78_c_fa1), .C(stage2_c78_c_fa2), .So(stage3_c79_s_fa0), .Co(stage3_c79_c_fa0));
    FA fa_1911(.A(stage2_c78_c_fa3), .B(stage2_c78_c_fa4), .C(stage2_c78_c_fa5), .So(stage3_c79_s_fa1), .Co(stage3_c79_c_fa1));
    FA fa_1912(.A(stage2_c78_c_fa6), .B(stage2_c78_c_fa7), .C(stage2_c79_s_fa0), .So(stage3_c79_s_fa2), .Co(stage3_c79_c_fa2));
    FA fa_1913(.A(stage2_c79_s_fa1), .B(stage2_c79_s_fa2), .C(stage2_c79_s_fa3), .So(stage3_c79_s_fa3), .Co(stage3_c79_c_fa3));
    FA fa_1914(.A(stage2_c79_s_fa4), .B(stage2_c79_s_fa5), .C(stage2_c79_s_fa6), .So(stage3_c79_s_fa4), .Co(stage3_c79_c_fa4));
    FA fa_1915(.A(stage2_c79_c_fa0), .B(stage2_c79_c_fa1), .C(stage2_c79_c_fa2), .So(stage3_c80_s_fa0), .Co(stage3_c80_c_fa0));
    FA fa_1916(.A(stage2_c79_c_fa3), .B(stage2_c79_c_fa4), .C(stage2_c79_c_fa5), .So(stage3_c80_s_fa1), .Co(stage3_c80_c_fa1));
    FA fa_1917(.A(stage2_c79_c_fa6), .B(stage2_c80_s_fa0), .C(stage2_c80_s_fa1), .So(stage3_c80_s_fa2), .Co(stage3_c80_c_fa2));
    FA fa_1918(.A(stage2_c80_s_fa2), .B(stage2_c80_s_fa3), .C(stage2_c80_s_fa4), .So(stage3_c80_s_fa3), .Co(stage3_c80_c_fa3));
    FA fa_1919(.A(stage2_c80_s_fa5), .B(stage2_c80_s_fa6), .C(stage1_c80_s_ha0), .So(stage3_c80_s_fa4), .Co(stage3_c80_c_fa4));
    FA fa_1920(.A(stage2_c80_c_fa0), .B(stage2_c80_c_fa1), .C(stage2_c80_c_fa2), .So(stage3_c81_s_fa0), .Co(stage3_c81_c_fa0));
    FA fa_1921(.A(stage2_c80_c_fa3), .B(stage2_c80_c_fa4), .C(stage2_c80_c_fa5), .So(stage3_c81_s_fa1), .Co(stage3_c81_c_fa1));
    FA fa_1922(.A(stage2_c80_c_fa6), .B(stage2_c81_s_fa0), .C(stage2_c81_s_fa1), .So(stage3_c81_s_fa2), .Co(stage3_c81_c_fa2));
    FA fa_1923(.A(stage2_c81_s_fa2), .B(stage2_c81_s_fa3), .C(stage2_c81_s_fa4), .So(stage3_c81_s_fa3), .Co(stage3_c81_c_fa3));
    FA fa_1924(.A(stage2_c81_s_fa5), .B(stage2_c81_s_fa6), .C(stage0_r71_c10), .So(stage3_c81_s_fa4), .Co(stage3_c81_c_fa4));
    FA fa_1925(.A(stage2_c81_c_fa0), .B(stage2_c81_c_fa1), .C(stage2_c81_c_fa2), .So(stage3_c82_s_fa0), .Co(stage3_c82_c_fa0));
    FA fa_1926(.A(stage2_c81_c_fa3), .B(stage2_c81_c_fa4), .C(stage2_c81_c_fa5), .So(stage3_c82_s_fa1), .Co(stage3_c82_c_fa1));
    FA fa_1927(.A(stage2_c81_c_fa6), .B(stage2_c82_s_fa0), .C(stage2_c82_s_fa1), .So(stage3_c82_s_fa2), .Co(stage3_c82_c_fa2));
    FA fa_1928(.A(stage2_c82_s_fa2), .B(stage2_c82_s_fa3), .C(stage2_c82_s_fa4), .So(stage3_c82_s_fa3), .Co(stage3_c82_c_fa3));
    HA ha_101(.A(stage2_c82_s_fa5), .B(stage2_c82_s_ha0), .So(stage3_c82_s_ha0), .Co(stage3_c82_c_ha0));
    FA fa_1929(.A(stage2_c82_c_fa0), .B(stage2_c82_c_fa1), .C(stage2_c82_c_fa2), .So(stage3_c83_s_fa0), .Co(stage3_c83_c_fa0));
    FA fa_1930(.A(stage2_c82_c_fa3), .B(stage2_c82_c_fa4), .C(stage2_c82_c_fa5), .So(stage3_c83_s_fa1), .Co(stage3_c83_c_fa1));
    FA fa_1931(.A(stage2_c82_c_ha0), .B(stage2_c83_s_fa0), .C(stage2_c83_s_fa1), .So(stage3_c83_s_fa2), .Co(stage3_c83_c_fa2));
    FA fa_1932(.A(stage2_c83_s_fa2), .B(stage2_c83_s_fa3), .C(stage2_c83_s_fa4), .So(stage3_c83_s_fa3), .Co(stage3_c83_c_fa3));
    HA ha_102(.A(stage2_c83_s_fa5), .B(stage2_c83_s_ha0), .So(stage3_c83_s_ha0), .Co(stage3_c83_c_ha0));
    FA fa_1933(.A(stage2_c83_c_fa0), .B(stage2_c83_c_fa1), .C(stage2_c83_c_fa2), .So(stage3_c84_s_fa0), .Co(stage3_c84_c_fa0));
    FA fa_1934(.A(stage2_c83_c_fa3), .B(stage2_c83_c_fa4), .C(stage2_c83_c_fa5), .So(stage3_c84_s_fa1), .Co(stage3_c84_c_fa1));
    FA fa_1935(.A(stage2_c83_c_ha0), .B(stage2_c84_s_fa0), .C(stage2_c84_s_fa1), .So(stage3_c84_s_fa2), .Co(stage3_c84_c_fa2));
    FA fa_1936(.A(stage2_c84_s_fa2), .B(stage2_c84_s_fa3), .C(stage2_c84_s_fa4), .So(stage3_c84_s_fa3), .Co(stage3_c84_c_fa3));
    HA ha_103(.A(stage2_c84_s_fa5), .B(stage2_c84_s_ha0), .So(stage3_c84_s_ha0), .Co(stage3_c84_c_ha0));
    FA fa_1937(.A(stage2_c84_c_fa0), .B(stage2_c84_c_fa1), .C(stage2_c84_c_fa2), .So(stage3_c85_s_fa0), .Co(stage3_c85_c_fa0));
    FA fa_1938(.A(stage2_c84_c_fa3), .B(stage2_c84_c_fa4), .C(stage2_c84_c_fa5), .So(stage3_c85_s_fa1), .Co(stage3_c85_c_fa1));
    FA fa_1939(.A(stage2_c84_c_ha0), .B(stage2_c85_s_fa0), .C(stage2_c85_s_fa1), .So(stage3_c85_s_fa2), .Co(stage3_c85_c_fa2));
    FA fa_1940(.A(stage2_c85_s_fa2), .B(stage2_c85_s_fa3), .C(stage2_c85_s_fa4), .So(stage3_c85_s_fa3), .Co(stage3_c85_c_fa3));
    FA fa_1941(.A(stage2_c85_c_fa0), .B(stage2_c85_c_fa1), .C(stage2_c85_c_fa2), .So(stage3_c86_s_fa0), .Co(stage3_c86_c_fa0));
    FA fa_1942(.A(stage2_c85_c_fa3), .B(stage2_c85_c_fa4), .C(stage2_c85_c_fa5), .So(stage3_c86_s_fa1), .Co(stage3_c86_c_fa1));
    FA fa_1943(.A(stage2_c86_s_fa0), .B(stage2_c86_s_fa1), .C(stage2_c86_s_fa2), .So(stage3_c86_s_fa2), .Co(stage3_c86_c_fa2));
    FA fa_1944(.A(stage2_c86_s_fa3), .B(stage2_c86_s_fa4), .C(stage2_c86_s_fa5), .So(stage3_c86_s_fa3), .Co(stage3_c86_c_fa3));
    FA fa_1945(.A(stage2_c86_c_fa0), .B(stage2_c86_c_fa1), .C(stage2_c86_c_fa2), .So(stage3_c87_s_fa0), .Co(stage3_c87_c_fa0));
    FA fa_1946(.A(stage2_c86_c_fa3), .B(stage2_c86_c_fa4), .C(stage2_c86_c_fa5), .So(stage3_c87_s_fa1), .Co(stage3_c87_c_fa1));
    FA fa_1947(.A(stage2_c87_s_fa0), .B(stage2_c87_s_fa1), .C(stage2_c87_s_fa2), .So(stage3_c87_s_fa2), .Co(stage3_c87_c_fa2));
    FA fa_1948(.A(stage2_c87_s_fa3), .B(stage2_c87_s_fa4), .C(stage2_c87_s_fa5), .So(stage3_c87_s_fa3), .Co(stage3_c87_c_fa3));
    FA fa_1949(.A(stage2_c87_c_fa0), .B(stage2_c87_c_fa1), .C(stage2_c87_c_fa2), .So(stage3_c88_s_fa0), .Co(stage3_c88_c_fa0));
    FA fa_1950(.A(stage2_c87_c_fa3), .B(stage2_c87_c_fa4), .C(stage2_c87_c_fa5), .So(stage3_c88_s_fa1), .Co(stage3_c88_c_fa1));
    FA fa_1951(.A(stage2_c88_s_fa0), .B(stage2_c88_s_fa1), .C(stage2_c88_s_fa2), .So(stage3_c88_s_fa2), .Co(stage3_c88_c_fa2));
    FA fa_1952(.A(stage2_c88_s_fa3), .B(stage2_c88_s_fa4), .C(stage1_c88_s_fa7), .So(stage3_c88_s_fa3), .Co(stage3_c88_c_fa3));
    FA fa_1953(.A(stage2_c88_c_fa0), .B(stage2_c88_c_fa1), .C(stage2_c88_c_fa2), .So(stage3_c89_s_fa0), .Co(stage3_c89_c_fa0));
    FA fa_1954(.A(stage2_c88_c_fa3), .B(stage2_c88_c_fa4), .C(stage2_c89_s_fa0), .So(stage3_c89_s_fa1), .Co(stage3_c89_c_fa1));
    FA fa_1955(.A(stage2_c89_s_fa1), .B(stage2_c89_s_fa2), .C(stage2_c89_s_fa3), .So(stage3_c89_s_fa2), .Co(stage3_c89_c_fa2));
    HA ha_104(.A(stage2_c89_s_fa4), .B(stage1_c89_s_ha0), .So(stage3_c89_s_ha0), .Co(stage3_c89_c_ha0));
    FA fa_1956(.A(stage2_c89_c_fa0), .B(stage2_c89_c_fa1), .C(stage2_c89_c_fa2), .So(stage3_c90_s_fa0), .Co(stage3_c90_c_fa0));
    FA fa_1957(.A(stage2_c89_c_fa3), .B(stage2_c89_c_fa4), .C(stage2_c90_s_fa0), .So(stage3_c90_s_fa1), .Co(stage3_c90_c_fa1));
    FA fa_1958(.A(stage2_c90_s_fa1), .B(stage2_c90_s_fa2), .C(stage2_c90_s_fa3), .So(stage3_c90_s_fa2), .Co(stage3_c90_c_fa2));
    HA ha_105(.A(stage2_c90_s_fa4), .B(stage0_r71_c19), .So(stage3_c90_s_ha0), .Co(stage3_c90_c_ha0));
    FA fa_1959(.A(stage2_c90_c_fa0), .B(stage2_c90_c_fa1), .C(stage2_c90_c_fa2), .So(stage3_c91_s_fa0), .Co(stage3_c91_c_fa0));
    FA fa_1960(.A(stage2_c90_c_fa3), .B(stage2_c90_c_fa4), .C(stage2_c91_s_fa0), .So(stage3_c91_s_fa1), .Co(stage3_c91_c_fa1));
    FA fa_1961(.A(stage2_c91_s_fa1), .B(stage2_c91_s_fa2), .C(stage2_c91_s_fa3), .So(stage3_c91_s_fa2), .Co(stage3_c91_c_fa2));
    FA fa_1962(.A(stage2_c91_c_fa0), .B(stage2_c91_c_fa1), .C(stage2_c91_c_fa2), .So(stage3_c92_s_fa0), .Co(stage3_c92_c_fa0));
    FA fa_1963(.A(stage2_c91_c_fa3), .B(stage2_c91_c_ha0), .C(stage2_c92_s_fa0), .So(stage3_c92_s_fa1), .Co(stage3_c92_c_fa1));
    FA fa_1964(.A(stage2_c92_s_fa1), .B(stage2_c92_s_fa2), .C(stage2_c92_s_fa3), .So(stage3_c92_s_fa2), .Co(stage3_c92_c_fa2));
    FA fa_1965(.A(stage2_c92_c_fa0), .B(stage2_c92_c_fa1), .C(stage2_c92_c_fa2), .So(stage3_c93_s_fa0), .Co(stage3_c93_c_fa0));
    FA fa_1966(.A(stage2_c92_c_fa3), .B(stage2_c92_c_ha0), .C(stage2_c93_s_fa0), .So(stage3_c93_s_fa1), .Co(stage3_c93_c_fa1));
    FA fa_1967(.A(stage2_c93_s_fa1), .B(stage2_c93_s_fa2), .C(stage2_c93_s_fa3), .So(stage3_c93_s_fa2), .Co(stage3_c93_c_fa2));
    FA fa_1968(.A(stage2_c93_c_fa0), .B(stage2_c93_c_fa1), .C(stage2_c93_c_fa2), .So(stage3_c94_s_fa0), .Co(stage3_c94_c_fa0));
    FA fa_1969(.A(stage2_c93_c_fa3), .B(stage2_c93_c_ha0), .C(stage2_c94_s_fa0), .So(stage3_c94_s_fa1), .Co(stage3_c94_c_fa1));
    FA fa_1970(.A(stage2_c94_s_fa1), .B(stage2_c94_s_fa2), .C(stage2_c94_s_fa3), .So(stage3_c94_s_fa2), .Co(stage3_c94_c_fa2));
    FA fa_1971(.A(stage2_c94_c_fa0), .B(stage2_c94_c_fa1), .C(stage2_c94_c_fa2), .So(stage3_c95_s_fa0), .Co(stage3_c95_c_fa0));
    FA fa_1972(.A(stage2_c94_c_fa3), .B(stage2_c95_s_fa0), .C(stage2_c95_s_fa1), .So(stage3_c95_s_fa1), .Co(stage3_c95_c_fa1));
    HA ha_106(.A(stage2_c95_s_fa2), .B(stage2_c95_s_fa3), .So(stage3_c95_s_ha0), .Co(stage3_c95_c_ha0));
    FA fa_1973(.A(stage2_c95_c_fa0), .B(stage2_c95_c_fa1), .C(stage2_c95_c_fa2), .So(stage3_c96_s_fa0), .Co(stage3_c96_c_fa0));
    FA fa_1974(.A(stage2_c95_c_fa3), .B(stage2_c96_s_fa0), .C(stage2_c96_s_fa1), .So(stage3_c96_s_fa1), .Co(stage3_c96_c_fa1));
    HA ha_107(.A(stage2_c96_s_fa2), .B(stage2_c96_s_fa3), .So(stage3_c96_s_ha0), .Co(stage3_c96_c_ha0));
    FA fa_1975(.A(stage2_c96_c_fa0), .B(stage2_c96_c_fa1), .C(stage2_c96_c_fa2), .So(stage3_c97_s_fa0), .Co(stage3_c97_c_fa0));
    FA fa_1976(.A(stage2_c96_c_fa3), .B(stage2_c97_s_fa0), .C(stage2_c97_s_fa1), .So(stage3_c97_s_fa1), .Co(stage3_c97_c_fa1));
    HA ha_108(.A(stage2_c97_s_fa2), .B(stage1_c97_s_fa4), .So(stage3_c97_s_ha0), .Co(stage3_c97_c_ha0));
    FA fa_1977(.A(stage2_c97_c_fa0), .B(stage2_c97_c_fa1), .C(stage2_c97_c_fa2), .So(stage3_c98_s_fa0), .Co(stage3_c98_c_fa0));
    FA fa_1978(.A(stage2_c98_s_fa0), .B(stage2_c98_s_fa1), .C(stage2_c98_s_fa2), .So(stage3_c98_s_fa1), .Co(stage3_c98_c_fa1));
    FA fa_1979(.A(stage2_c98_c_fa0), .B(stage2_c98_c_fa1), .C(stage2_c98_c_fa2), .So(stage3_c99_s_fa0), .Co(stage3_c99_c_fa0));
    FA fa_1980(.A(stage2_c99_s_fa0), .B(stage2_c99_s_fa1), .C(stage2_c99_s_fa2), .So(stage3_c99_s_fa1), .Co(stage3_c99_c_fa1));
    FA fa_1981(.A(stage2_c99_c_fa0), .B(stage2_c99_c_fa1), .C(stage2_c99_c_fa2), .So(stage3_c100_s_fa0), .Co(stage3_c100_c_fa0));
    FA fa_1982(.A(stage2_c100_s_fa0), .B(stage2_c100_s_fa1), .C(stage2_c100_s_ha0), .So(stage3_c100_s_fa1), .Co(stage3_c100_c_fa1));
    FA fa_1983(.A(stage2_c100_c_fa0), .B(stage2_c100_c_fa1), .C(stage2_c100_c_ha0), .So(stage3_c101_s_fa0), .Co(stage3_c101_c_fa0));
    FA fa_1984(.A(stage2_c101_s_fa0), .B(stage2_c101_s_fa1), .C(stage2_c101_s_ha0), .So(stage3_c101_s_fa1), .Co(stage3_c101_c_fa1));
    FA fa_1985(.A(stage2_c101_c_fa0), .B(stage2_c101_c_fa1), .C(stage2_c101_c_ha0), .So(stage3_c102_s_fa0), .Co(stage3_c102_c_fa0));
    FA fa_1986(.A(stage2_c102_s_fa0), .B(stage2_c102_s_fa1), .C(stage2_c102_s_ha0), .So(stage3_c102_s_fa1), .Co(stage3_c102_c_fa1));
    FA fa_1987(.A(stage2_c102_c_fa0), .B(stage2_c102_c_fa1), .C(stage2_c102_c_ha0), .So(stage3_c103_s_fa0), .Co(stage3_c103_c_fa0));
    HA ha_109(.A(stage2_c103_s_fa0), .B(stage2_c103_s_fa1), .So(stage3_c103_s_ha0), .Co(stage3_c103_c_ha0));
    FA fa_1988(.A(stage2_c103_c_fa0), .B(stage2_c103_c_fa1), .C(stage2_c104_s_fa0), .So(stage3_c104_s_fa0), .Co(stage3_c104_c_fa0));
    FA fa_1989(.A(stage2_c104_c_fa0), .B(stage2_c104_c_fa1), .C(stage2_c105_s_fa0), .So(stage3_c105_s_fa0), .Co(stage3_c105_c_fa0));
    FA fa_1990(.A(stage2_c105_c_fa0), .B(stage2_c105_c_fa1), .C(stage2_c106_s_fa0), .So(stage3_c106_s_fa0), .Co(stage3_c106_c_fa0));
    FA fa_1991(.A(stage2_c106_c_fa0), .B(stage2_c107_s_fa0), .C(stage1_c107_s_ha0), .So(stage3_c107_s_fa0), .Co(stage3_c107_c_fa0));
    FA fa_1992(.A(stage2_c107_c_fa0), .B(stage2_c108_s_fa0), .C(stage0_r71_c37), .So(stage3_c108_s_fa0), .Co(stage3_c108_c_fa0));
    HA ha_110(.A(stage2_c108_c_fa0), .B(stage2_c109_s_ha0), .So(stage3_c109_s_ha0), .Co(stage3_c109_c_ha0));
    HA ha_111(.A(stage2_c109_c_ha0), .B(stage2_c110_s_ha0), .So(stage3_c110_s_ha0), .Co(stage3_c110_c_ha0));
    HA ha_112(.A(stage2_c110_c_ha0), .B(stage2_c111_s_ha0), .So(stage3_c111_s_ha0), .Co(stage3_c111_c_ha0));
    HA ha_113(.A(stage3_c3_c_ha0), .B(stage3_c4_s_ha0), .So(stage4_c4_s_ha0), .Co(stage4_c4_c_ha0));
    HA ha_114(.A(stage3_c4_c_ha0), .B(stage3_c5_s_fa0), .So(stage4_c5_s_ha0), .Co(stage4_c5_c_ha0));
    HA ha_115(.A(stage3_c5_c_fa0), .B(stage3_c6_s_fa0), .So(stage4_c6_s_ha0), .Co(stage4_c6_c_ha0));
    FA fa_1993(.A(stage3_c6_c_fa0), .B(stage3_c7_s_fa0), .C(stage2_c7_s_ha0), .So(stage4_c7_s_fa0), .Co(stage4_c7_c_fa0));
    FA fa_1994(.A(stage3_c7_c_fa0), .B(stage3_c8_s_fa0), .C(stage2_c8_s_fa1), .So(stage4_c8_s_fa0), .Co(stage4_c8_c_fa0));
    FA fa_1995(.A(stage3_c8_c_fa0), .B(stage3_c9_s_fa0), .C(stage3_c9_s_ha0), .So(stage4_c9_s_fa0), .Co(stage4_c9_c_fa0));
    FA fa_1996(.A(stage3_c9_c_fa0), .B(stage3_c9_c_ha0), .C(stage3_c10_s_fa0), .So(stage4_c10_s_fa0), .Co(stage4_c10_c_fa0));
    FA fa_1997(.A(stage3_c10_c_fa0), .B(stage3_c10_c_ha0), .C(stage3_c11_s_fa0), .So(stage4_c11_s_fa0), .Co(stage4_c11_c_fa0));
    FA fa_1998(.A(stage3_c11_c_fa0), .B(stage3_c11_c_ha0), .C(stage3_c12_s_fa0), .So(stage4_c12_s_fa0), .Co(stage4_c12_c_fa0));
    FA fa_1999(.A(stage3_c12_c_fa0), .B(stage3_c12_c_fa1), .C(stage3_c13_s_fa0), .So(stage4_c13_s_fa0), .Co(stage4_c13_c_fa0));
    FA fa_2000(.A(stage3_c13_c_fa0), .B(stage3_c13_c_fa1), .C(stage3_c14_s_fa0), .So(stage4_c14_s_fa0), .Co(stage4_c14_c_fa0));
    HA ha_116(.A(stage3_c14_s_fa1), .B(stage1_c14_s_fa4), .So(stage4_c14_s_ha0), .Co(stage4_c14_c_ha0));
    FA fa_2001(.A(stage3_c14_c_fa0), .B(stage3_c14_c_fa1), .C(stage3_c15_s_fa0), .So(stage4_c15_s_fa0), .Co(stage4_c15_c_fa0));
    HA ha_117(.A(stage3_c15_s_fa1), .B(stage2_c15_s_ha0), .So(stage4_c15_s_ha0), .Co(stage4_c15_c_ha0));
    FA fa_2002(.A(stage3_c15_c_fa0), .B(stage3_c15_c_fa1), .C(stage3_c16_s_fa0), .So(stage4_c16_s_fa0), .Co(stage4_c16_c_fa0));
    HA ha_118(.A(stage3_c16_s_fa1), .B(stage3_c16_s_ha0), .So(stage4_c16_s_ha0), .Co(stage4_c16_c_ha0));
    FA fa_2003(.A(stage3_c16_c_fa0), .B(stage3_c16_c_fa1), .C(stage3_c16_c_ha0), .So(stage4_c17_s_fa0), .Co(stage4_c17_c_fa0));
    FA fa_2004(.A(stage3_c17_s_fa0), .B(stage3_c17_s_fa1), .C(stage3_c17_s_ha0), .So(stage4_c17_s_fa1), .Co(stage4_c17_c_fa1));
    FA fa_2005(.A(stage3_c17_c_fa0), .B(stage3_c17_c_fa1), .C(stage3_c17_c_ha0), .So(stage4_c18_s_fa0), .Co(stage4_c18_c_fa0));
    FA fa_2006(.A(stage3_c18_s_fa0), .B(stage3_c18_s_fa1), .C(stage3_c18_s_fa2), .So(stage4_c18_s_fa1), .Co(stage4_c18_c_fa1));
    FA fa_2007(.A(stage3_c18_c_fa0), .B(stage3_c18_c_fa1), .C(stage3_c18_c_fa2), .So(stage4_c19_s_fa0), .Co(stage4_c19_c_fa0));
    FA fa_2008(.A(stage3_c19_s_fa0), .B(stage3_c19_s_fa1), .C(stage3_c19_s_fa2), .So(stage4_c19_s_fa1), .Co(stage4_c19_c_fa1));
    FA fa_2009(.A(stage3_c19_c_fa0), .B(stage3_c19_c_fa1), .C(stage3_c19_c_fa2), .So(stage4_c20_s_fa0), .Co(stage4_c20_c_fa0));
    FA fa_2010(.A(stage3_c20_s_fa0), .B(stage3_c20_s_fa1), .C(stage3_c20_s_fa2), .So(stage4_c20_s_fa1), .Co(stage4_c20_c_fa1));
    FA fa_2011(.A(stage3_c20_c_fa0), .B(stage3_c20_c_fa1), .C(stage3_c20_c_fa2), .So(stage4_c21_s_fa0), .Co(stage4_c21_c_fa0));
    FA fa_2012(.A(stage3_c21_s_fa0), .B(stage3_c21_s_fa1), .C(stage3_c21_s_fa2), .So(stage4_c21_s_fa1), .Co(stage4_c21_c_fa1));
    FA fa_2013(.A(stage3_c21_c_fa0), .B(stage3_c21_c_fa1), .C(stage3_c21_c_fa2), .So(stage4_c22_s_fa0), .Co(stage4_c22_c_fa0));
    FA fa_2014(.A(stage3_c22_s_fa0), .B(stage3_c22_s_fa1), .C(stage3_c22_s_fa2), .So(stage4_c22_s_fa1), .Co(stage4_c22_c_fa1));
    FA fa_2015(.A(stage3_c22_c_fa0), .B(stage3_c22_c_fa1), .C(stage3_c22_c_fa2), .So(stage4_c23_s_fa0), .Co(stage4_c23_c_fa0));
    FA fa_2016(.A(stage3_c23_s_fa0), .B(stage3_c23_s_fa1), .C(stage3_c23_s_fa2), .So(stage4_c23_s_fa1), .Co(stage4_c23_c_fa1));
    FA fa_2017(.A(stage3_c23_c_fa0), .B(stage3_c23_c_fa1), .C(stage3_c23_c_fa2), .So(stage4_c24_s_fa0), .Co(stage4_c24_c_fa0));
    FA fa_2018(.A(stage3_c23_c_ha0), .B(stage3_c24_s_fa0), .C(stage3_c24_s_fa1), .So(stage4_c24_s_fa1), .Co(stage4_c24_c_fa1));
    HA ha_119(.A(stage3_c24_s_fa2), .B(stage3_c24_s_ha0), .So(stage4_c24_s_ha0), .Co(stage4_c24_c_ha0));
    FA fa_2019(.A(stage3_c24_c_fa0), .B(stage3_c24_c_fa1), .C(stage3_c24_c_fa2), .So(stage4_c25_s_fa0), .Co(stage4_c25_c_fa0));
    FA fa_2020(.A(stage3_c24_c_ha0), .B(stage3_c25_s_fa0), .C(stage3_c25_s_fa1), .So(stage4_c25_s_fa1), .Co(stage4_c25_c_fa1));
    HA ha_120(.A(stage3_c25_s_fa2), .B(stage3_c25_s_fa3), .So(stage4_c25_s_ha0), .Co(stage4_c25_c_ha0));
    FA fa_2021(.A(stage3_c25_c_fa0), .B(stage3_c25_c_fa1), .C(stage3_c25_c_fa2), .So(stage4_c26_s_fa0), .Co(stage4_c26_c_fa0));
    FA fa_2022(.A(stage3_c25_c_fa3), .B(stage3_c26_s_fa0), .C(stage3_c26_s_fa1), .So(stage4_c26_s_fa1), .Co(stage4_c26_c_fa1));
    HA ha_121(.A(stage3_c26_s_fa2), .B(stage3_c26_s_fa3), .So(stage4_c26_s_ha0), .Co(stage4_c26_c_ha0));
    FA fa_2023(.A(stage3_c26_c_fa0), .B(stage3_c26_c_fa1), .C(stage3_c26_c_fa2), .So(stage4_c27_s_fa0), .Co(stage4_c27_c_fa0));
    FA fa_2024(.A(stage3_c26_c_fa3), .B(stage3_c27_s_fa0), .C(stage3_c27_s_fa1), .So(stage4_c27_s_fa1), .Co(stage4_c27_c_fa1));
    FA fa_2025(.A(stage3_c27_s_fa2), .B(stage3_c27_s_fa3), .C(stage0_r27_c0), .So(stage4_c27_s_fa2), .Co(stage4_c27_c_fa2));
    FA fa_2026(.A(stage3_c27_c_fa0), .B(stage3_c27_c_fa1), .C(stage3_c27_c_fa2), .So(stage4_c28_s_fa0), .Co(stage4_c28_c_fa0));
    FA fa_2027(.A(stage3_c27_c_fa3), .B(stage3_c28_s_fa0), .C(stage3_c28_s_fa1), .So(stage4_c28_s_fa1), .Co(stage4_c28_c_fa1));
    FA fa_2028(.A(stage3_c28_s_fa2), .B(stage3_c28_s_fa3), .C(stage1_c28_s_ha0), .So(stage4_c28_s_fa2), .Co(stage4_c28_c_fa2));
    FA fa_2029(.A(stage3_c28_c_fa0), .B(stage3_c28_c_fa1), .C(stage3_c28_c_fa2), .So(stage4_c29_s_fa0), .Co(stage4_c29_c_fa0));
    FA fa_2030(.A(stage3_c28_c_fa3), .B(stage3_c29_s_fa0), .C(stage3_c29_s_fa1), .So(stage4_c29_s_fa1), .Co(stage4_c29_c_fa1));
    FA fa_2031(.A(stage3_c29_s_fa2), .B(stage3_c29_s_fa3), .C(stage2_c29_s_ha0), .So(stage4_c29_s_fa2), .Co(stage4_c29_c_fa2));
    FA fa_2032(.A(stage3_c29_c_fa0), .B(stage3_c29_c_fa1), .C(stage3_c29_c_fa2), .So(stage4_c30_s_fa0), .Co(stage4_c30_c_fa0));
    FA fa_2033(.A(stage3_c29_c_fa3), .B(stage3_c30_s_fa0), .C(stage3_c30_s_fa1), .So(stage4_c30_s_fa1), .Co(stage4_c30_c_fa1));
    FA fa_2034(.A(stage3_c30_s_fa2), .B(stage3_c30_s_fa3), .C(stage3_c30_s_ha0), .So(stage4_c30_s_fa2), .Co(stage4_c30_c_fa2));
    FA fa_2035(.A(stage3_c30_c_fa0), .B(stage3_c30_c_fa1), .C(stage3_c30_c_fa2), .So(stage4_c31_s_fa0), .Co(stage4_c31_c_fa0));
    FA fa_2036(.A(stage3_c30_c_fa3), .B(stage3_c30_c_ha0), .C(stage3_c31_s_fa0), .So(stage4_c31_s_fa1), .Co(stage4_c31_c_fa1));
    FA fa_2037(.A(stage3_c31_s_fa1), .B(stage3_c31_s_fa2), .C(stage3_c31_s_fa3), .So(stage4_c31_s_fa2), .Co(stage4_c31_c_fa2));
    FA fa_2038(.A(stage3_c31_c_fa0), .B(stage3_c31_c_fa1), .C(stage3_c31_c_fa2), .So(stage4_c32_s_fa0), .Co(stage4_c32_c_fa0));
    FA fa_2039(.A(stage3_c31_c_fa3), .B(stage3_c31_c_ha0), .C(stage3_c32_s_fa0), .So(stage4_c32_s_fa1), .Co(stage4_c32_c_fa1));
    FA fa_2040(.A(stage3_c32_s_fa1), .B(stage3_c32_s_fa2), .C(stage3_c32_s_fa3), .So(stage4_c32_s_fa2), .Co(stage4_c32_c_fa2));
    FA fa_2041(.A(stage3_c32_c_fa0), .B(stage3_c32_c_fa1), .C(stage3_c32_c_fa2), .So(stage4_c33_s_fa0), .Co(stage4_c33_c_fa0));
    FA fa_2042(.A(stage3_c32_c_fa3), .B(stage3_c32_c_fa4), .C(stage3_c33_s_fa0), .So(stage4_c33_s_fa1), .Co(stage4_c33_c_fa1));
    FA fa_2043(.A(stage3_c33_s_fa1), .B(stage3_c33_s_fa2), .C(stage3_c33_s_fa3), .So(stage4_c33_s_fa2), .Co(stage4_c33_c_fa2));
    FA fa_2044(.A(stage3_c33_c_fa0), .B(stage3_c33_c_fa1), .C(stage3_c33_c_fa2), .So(stage4_c34_s_fa0), .Co(stage4_c34_c_fa0));
    FA fa_2045(.A(stage3_c33_c_fa3), .B(stage3_c33_c_fa4), .C(stage3_c34_s_fa0), .So(stage4_c34_s_fa1), .Co(stage4_c34_c_fa1));
    FA fa_2046(.A(stage3_c34_s_fa1), .B(stage3_c34_s_fa2), .C(stage3_c34_s_fa3), .So(stage4_c34_s_fa2), .Co(stage4_c34_c_fa2));
    HA ha_122(.A(stage3_c34_s_fa4), .B(stage2_c34_s_ha0), .So(stage4_c34_s_ha0), .Co(stage4_c34_c_ha0));
    FA fa_2047(.A(stage3_c34_c_fa0), .B(stage3_c34_c_fa1), .C(stage3_c34_c_fa2), .So(stage4_c35_s_fa0), .Co(stage4_c35_c_fa0));
    FA fa_2048(.A(stage3_c34_c_fa3), .B(stage3_c34_c_fa4), .C(stage3_c35_s_fa0), .So(stage4_c35_s_fa1), .Co(stage4_c35_c_fa1));
    FA fa_2049(.A(stage3_c35_s_fa1), .B(stage3_c35_s_fa2), .C(stage3_c35_s_fa3), .So(stage4_c35_s_fa2), .Co(stage4_c35_c_fa2));
    HA ha_123(.A(stage3_c35_s_fa4), .B(stage2_c35_s_fa7), .So(stage4_c35_s_ha0), .Co(stage4_c35_c_ha0));
    FA fa_2050(.A(stage3_c35_c_fa0), .B(stage3_c35_c_fa1), .C(stage3_c35_c_fa2), .So(stage4_c36_s_fa0), .Co(stage4_c36_c_fa0));
    FA fa_2051(.A(stage3_c35_c_fa3), .B(stage3_c35_c_fa4), .C(stage3_c36_s_fa0), .So(stage4_c36_s_fa1), .Co(stage4_c36_c_fa1));
    FA fa_2052(.A(stage3_c36_s_fa1), .B(stage3_c36_s_fa2), .C(stage3_c36_s_fa3), .So(stage4_c36_s_fa2), .Co(stage4_c36_c_fa2));
    HA ha_124(.A(stage3_c36_s_fa4), .B(stage3_c36_s_ha0), .So(stage4_c36_s_ha0), .Co(stage4_c36_c_ha0));
    FA fa_2053(.A(stage3_c36_c_fa0), .B(stage3_c36_c_fa1), .C(stage3_c36_c_fa2), .So(stage4_c37_s_fa0), .Co(stage4_c37_c_fa0));
    FA fa_2054(.A(stage3_c36_c_fa3), .B(stage3_c36_c_fa4), .C(stage3_c36_c_ha0), .So(stage4_c37_s_fa1), .Co(stage4_c37_c_fa1));
    FA fa_2055(.A(stage3_c37_s_fa0), .B(stage3_c37_s_fa1), .C(stage3_c37_s_fa2), .So(stage4_c37_s_fa2), .Co(stage4_c37_c_fa2));
    FA fa_2056(.A(stage3_c37_s_fa3), .B(stage3_c37_s_fa4), .C(stage3_c37_s_ha0), .So(stage4_c37_s_fa3), .Co(stage4_c37_c_fa3));
    FA fa_2057(.A(stage3_c37_c_fa0), .B(stage3_c37_c_fa1), .C(stage3_c37_c_fa2), .So(stage4_c38_s_fa0), .Co(stage4_c38_c_fa0));
    FA fa_2058(.A(stage3_c37_c_fa3), .B(stage3_c37_c_fa4), .C(stage3_c37_c_ha0), .So(stage4_c38_s_fa1), .Co(stage4_c38_c_fa1));
    FA fa_2059(.A(stage3_c38_s_fa0), .B(stage3_c38_s_fa1), .C(stage3_c38_s_fa2), .So(stage4_c38_s_fa2), .Co(stage4_c38_c_fa2));
    FA fa_2060(.A(stage3_c38_s_fa3), .B(stage3_c38_s_fa4), .C(stage3_c38_s_ha0), .So(stage4_c38_s_fa3), .Co(stage4_c38_c_fa3));
    FA fa_2061(.A(stage3_c38_c_fa0), .B(stage3_c38_c_fa1), .C(stage3_c38_c_fa2), .So(stage4_c39_s_fa0), .Co(stage4_c39_c_fa0));
    FA fa_2062(.A(stage3_c38_c_fa3), .B(stage3_c38_c_fa4), .C(stage3_c38_c_ha0), .So(stage4_c39_s_fa1), .Co(stage4_c39_c_fa1));
    FA fa_2063(.A(stage3_c39_s_fa0), .B(stage3_c39_s_fa1), .C(stage3_c39_s_fa2), .So(stage4_c39_s_fa2), .Co(stage4_c39_c_fa2));
    FA fa_2064(.A(stage3_c39_s_fa3), .B(stage3_c39_s_fa4), .C(stage3_c39_s_fa5), .So(stage4_c39_s_fa3), .Co(stage4_c39_c_fa3));
    FA fa_2065(.A(stage3_c39_c_fa0), .B(stage3_c39_c_fa1), .C(stage3_c39_c_fa2), .So(stage4_c40_s_fa0), .Co(stage4_c40_c_fa0));
    FA fa_2066(.A(stage3_c39_c_fa3), .B(stage3_c39_c_fa4), .C(stage3_c39_c_fa5), .So(stage4_c40_s_fa1), .Co(stage4_c40_c_fa1));
    FA fa_2067(.A(stage3_c40_s_fa0), .B(stage3_c40_s_fa1), .C(stage3_c40_s_fa2), .So(stage4_c40_s_fa2), .Co(stage4_c40_c_fa2));
    FA fa_2068(.A(stage3_c40_s_fa3), .B(stage3_c40_s_fa4), .C(stage3_c40_s_fa5), .So(stage4_c40_s_fa3), .Co(stage4_c40_c_fa3));
    FA fa_2069(.A(stage3_c40_c_fa0), .B(stage3_c40_c_fa1), .C(stage3_c40_c_fa2), .So(stage4_c41_s_fa0), .Co(stage4_c41_c_fa0));
    FA fa_2070(.A(stage3_c40_c_fa3), .B(stage3_c40_c_fa4), .C(stage3_c40_c_fa5), .So(stage4_c41_s_fa1), .Co(stage4_c41_c_fa1));
    FA fa_2071(.A(stage3_c41_s_fa0), .B(stage3_c41_s_fa1), .C(stage3_c41_s_fa2), .So(stage4_c41_s_fa2), .Co(stage4_c41_c_fa2));
    FA fa_2072(.A(stage3_c41_s_fa3), .B(stage3_c41_s_fa4), .C(stage3_c41_s_fa5), .So(stage4_c41_s_fa3), .Co(stage4_c41_c_fa3));
    FA fa_2073(.A(stage3_c41_c_fa0), .B(stage3_c41_c_fa1), .C(stage3_c41_c_fa2), .So(stage4_c42_s_fa0), .Co(stage4_c42_c_fa0));
    FA fa_2074(.A(stage3_c41_c_fa3), .B(stage3_c41_c_fa4), .C(stage3_c41_c_fa5), .So(stage4_c42_s_fa1), .Co(stage4_c42_c_fa1));
    FA fa_2075(.A(stage3_c42_s_fa0), .B(stage3_c42_s_fa1), .C(stage3_c42_s_fa2), .So(stage4_c42_s_fa2), .Co(stage4_c42_c_fa2));
    FA fa_2076(.A(stage3_c42_s_fa3), .B(stage3_c42_s_fa4), .C(stage3_c42_s_fa5), .So(stage4_c42_s_fa3), .Co(stage4_c42_c_fa3));
    FA fa_2077(.A(stage3_c42_c_fa0), .B(stage3_c42_c_fa1), .C(stage3_c42_c_fa2), .So(stage4_c43_s_fa0), .Co(stage4_c43_c_fa0));
    FA fa_2078(.A(stage3_c42_c_fa3), .B(stage3_c42_c_fa4), .C(stage3_c42_c_fa5), .So(stage4_c43_s_fa1), .Co(stage4_c43_c_fa1));
    FA fa_2079(.A(stage3_c43_s_fa0), .B(stage3_c43_s_fa1), .C(stage3_c43_s_fa2), .So(stage4_c43_s_fa2), .Co(stage4_c43_c_fa2));
    FA fa_2080(.A(stage3_c43_s_fa3), .B(stage3_c43_s_fa4), .C(stage3_c43_s_fa5), .So(stage4_c43_s_fa3), .Co(stage4_c43_c_fa3));
    FA fa_2081(.A(stage3_c43_c_fa0), .B(stage3_c43_c_fa1), .C(stage3_c43_c_fa2), .So(stage4_c44_s_fa0), .Co(stage4_c44_c_fa0));
    FA fa_2082(.A(stage3_c43_c_fa3), .B(stage3_c43_c_fa4), .C(stage3_c43_c_fa5), .So(stage4_c44_s_fa1), .Co(stage4_c44_c_fa1));
    FA fa_2083(.A(stage3_c44_s_fa0), .B(stage3_c44_s_fa1), .C(stage3_c44_s_fa2), .So(stage4_c44_s_fa2), .Co(stage4_c44_c_fa2));
    FA fa_2084(.A(stage3_c44_s_fa3), .B(stage3_c44_s_fa4), .C(stage3_c44_s_fa5), .So(stage4_c44_s_fa3), .Co(stage4_c44_c_fa3));
    FA fa_2085(.A(stage3_c44_c_fa0), .B(stage3_c44_c_fa1), .C(stage3_c44_c_fa2), .So(stage4_c45_s_fa0), .Co(stage4_c45_c_fa0));
    FA fa_2086(.A(stage3_c44_c_fa3), .B(stage3_c44_c_fa4), .C(stage3_c44_c_fa5), .So(stage4_c45_s_fa1), .Co(stage4_c45_c_fa1));
    FA fa_2087(.A(stage3_c45_s_fa0), .B(stage3_c45_s_fa1), .C(stage3_c45_s_fa2), .So(stage4_c45_s_fa2), .Co(stage4_c45_c_fa2));
    FA fa_2088(.A(stage3_c45_s_fa3), .B(stage3_c45_s_fa4), .C(stage3_c45_s_fa5), .So(stage4_c45_s_fa3), .Co(stage4_c45_c_fa3));
    FA fa_2089(.A(stage3_c45_c_fa0), .B(stage3_c45_c_fa1), .C(stage3_c45_c_fa2), .So(stage4_c46_s_fa0), .Co(stage4_c46_c_fa0));
    FA fa_2090(.A(stage3_c45_c_fa3), .B(stage3_c45_c_fa4), .C(stage3_c45_c_fa5), .So(stage4_c46_s_fa1), .Co(stage4_c46_c_fa1));
    FA fa_2091(.A(stage3_c46_s_fa0), .B(stage3_c46_s_fa1), .C(stage3_c46_s_fa2), .So(stage4_c46_s_fa2), .Co(stage4_c46_c_fa2));
    FA fa_2092(.A(stage3_c46_s_fa3), .B(stage3_c46_s_fa4), .C(stage3_c46_s_fa5), .So(stage4_c46_s_fa3), .Co(stage4_c46_c_fa3));
    FA fa_2093(.A(stage3_c46_c_fa0), .B(stage3_c46_c_fa1), .C(stage3_c46_c_fa2), .So(stage4_c47_s_fa0), .Co(stage4_c47_c_fa0));
    FA fa_2094(.A(stage3_c46_c_fa3), .B(stage3_c46_c_fa4), .C(stage3_c46_c_fa5), .So(stage4_c47_s_fa1), .Co(stage4_c47_c_fa1));
    FA fa_2095(.A(stage3_c47_s_fa0), .B(stage3_c47_s_fa1), .C(stage3_c47_s_fa2), .So(stage4_c47_s_fa2), .Co(stage4_c47_c_fa2));
    FA fa_2096(.A(stage3_c47_s_fa3), .B(stage3_c47_s_fa4), .C(stage3_c47_s_fa5), .So(stage4_c47_s_fa3), .Co(stage4_c47_c_fa3));
    FA fa_2097(.A(stage3_c47_c_fa0), .B(stage3_c47_c_fa1), .C(stage3_c47_c_fa2), .So(stage4_c48_s_fa0), .Co(stage4_c48_c_fa0));
    FA fa_2098(.A(stage3_c47_c_fa3), .B(stage3_c47_c_fa4), .C(stage3_c47_c_fa5), .So(stage4_c48_s_fa1), .Co(stage4_c48_c_fa1));
    FA fa_2099(.A(stage3_c48_s_fa0), .B(stage3_c48_s_fa1), .C(stage3_c48_s_fa2), .So(stage4_c48_s_fa2), .Co(stage4_c48_c_fa2));
    FA fa_2100(.A(stage3_c48_s_fa3), .B(stage3_c48_s_fa4), .C(stage3_c48_s_fa5), .So(stage4_c48_s_fa3), .Co(stage4_c48_c_fa3));
    FA fa_2101(.A(stage3_c48_c_fa0), .B(stage3_c48_c_fa1), .C(stage3_c48_c_fa2), .So(stage4_c49_s_fa0), .Co(stage4_c49_c_fa0));
    FA fa_2102(.A(stage3_c48_c_fa3), .B(stage3_c48_c_fa4), .C(stage3_c48_c_fa5), .So(stage4_c49_s_fa1), .Co(stage4_c49_c_fa1));
    FA fa_2103(.A(stage3_c49_s_fa0), .B(stage3_c49_s_fa1), .C(stage3_c49_s_fa2), .So(stage4_c49_s_fa2), .Co(stage4_c49_c_fa2));
    FA fa_2104(.A(stage3_c49_s_fa3), .B(stage3_c49_s_fa4), .C(stage3_c49_s_fa5), .So(stage4_c49_s_fa3), .Co(stage4_c49_c_fa3));
    FA fa_2105(.A(stage3_c49_c_fa0), .B(stage3_c49_c_fa1), .C(stage3_c49_c_fa2), .So(stage4_c50_s_fa0), .Co(stage4_c50_c_fa0));
    FA fa_2106(.A(stage3_c49_c_fa3), .B(stage3_c49_c_fa4), .C(stage3_c49_c_fa5), .So(stage4_c50_s_fa1), .Co(stage4_c50_c_fa1));
    FA fa_2107(.A(stage3_c50_s_fa0), .B(stage3_c50_s_fa1), .C(stage3_c50_s_fa2), .So(stage4_c50_s_fa2), .Co(stage4_c50_c_fa2));
    FA fa_2108(.A(stage3_c50_s_fa3), .B(stage3_c50_s_fa4), .C(stage3_c50_s_fa5), .So(stage4_c50_s_fa3), .Co(stage4_c50_c_fa3));
    FA fa_2109(.A(stage3_c50_c_fa0), .B(stage3_c50_c_fa1), .C(stage3_c50_c_fa2), .So(stage4_c51_s_fa0), .Co(stage4_c51_c_fa0));
    FA fa_2110(.A(stage3_c50_c_fa3), .B(stage3_c50_c_fa4), .C(stage3_c50_c_fa5), .So(stage4_c51_s_fa1), .Co(stage4_c51_c_fa1));
    FA fa_2111(.A(stage3_c51_s_fa0), .B(stage3_c51_s_fa1), .C(stage3_c51_s_fa2), .So(stage4_c51_s_fa2), .Co(stage4_c51_c_fa2));
    FA fa_2112(.A(stage3_c51_s_fa3), .B(stage3_c51_s_fa4), .C(stage3_c51_s_fa5), .So(stage4_c51_s_fa3), .Co(stage4_c51_c_fa3));
    FA fa_2113(.A(stage3_c51_c_fa0), .B(stage3_c51_c_fa1), .C(stage3_c51_c_fa2), .So(stage4_c52_s_fa0), .Co(stage4_c52_c_fa0));
    FA fa_2114(.A(stage3_c51_c_fa3), .B(stage3_c51_c_fa4), .C(stage3_c51_c_fa5), .So(stage4_c52_s_fa1), .Co(stage4_c52_c_fa1));
    FA fa_2115(.A(stage3_c52_s_fa0), .B(stage3_c52_s_fa1), .C(stage3_c52_s_fa2), .So(stage4_c52_s_fa2), .Co(stage4_c52_c_fa2));
    FA fa_2116(.A(stage3_c52_s_fa3), .B(stage3_c52_s_fa4), .C(stage3_c52_s_fa5), .So(stage4_c52_s_fa3), .Co(stage4_c52_c_fa3));
    FA fa_2117(.A(stage3_c52_c_fa0), .B(stage3_c52_c_fa1), .C(stage3_c52_c_fa2), .So(stage4_c53_s_fa0), .Co(stage4_c53_c_fa0));
    FA fa_2118(.A(stage3_c52_c_fa3), .B(stage3_c52_c_fa4), .C(stage3_c52_c_fa5), .So(stage4_c53_s_fa1), .Co(stage4_c53_c_fa1));
    FA fa_2119(.A(stage3_c53_s_fa0), .B(stage3_c53_s_fa1), .C(stage3_c53_s_fa2), .So(stage4_c53_s_fa2), .Co(stage4_c53_c_fa2));
    FA fa_2120(.A(stage3_c53_s_fa3), .B(stage3_c53_s_fa4), .C(stage3_c53_s_fa5), .So(stage4_c53_s_fa3), .Co(stage4_c53_c_fa3));
    FA fa_2121(.A(stage3_c53_c_fa0), .B(stage3_c53_c_fa1), .C(stage3_c53_c_fa2), .So(stage4_c54_s_fa0), .Co(stage4_c54_c_fa0));
    FA fa_2122(.A(stage3_c53_c_fa3), .B(stage3_c53_c_fa4), .C(stage3_c53_c_fa5), .So(stage4_c54_s_fa1), .Co(stage4_c54_c_fa1));
    FA fa_2123(.A(stage3_c54_s_fa0), .B(stage3_c54_s_fa1), .C(stage3_c54_s_fa2), .So(stage4_c54_s_fa2), .Co(stage4_c54_c_fa2));
    FA fa_2124(.A(stage3_c54_s_fa3), .B(stage3_c54_s_fa4), .C(stage3_c54_s_fa5), .So(stage4_c54_s_fa3), .Co(stage4_c54_c_fa3));
    FA fa_2125(.A(stage3_c54_c_fa0), .B(stage3_c54_c_fa1), .C(stage3_c54_c_fa2), .So(stage4_c55_s_fa0), .Co(stage4_c55_c_fa0));
    FA fa_2126(.A(stage3_c54_c_fa3), .B(stage3_c54_c_fa4), .C(stage3_c54_c_fa5), .So(stage4_c55_s_fa1), .Co(stage4_c55_c_fa1));
    FA fa_2127(.A(stage3_c55_s_fa0), .B(stage3_c55_s_fa1), .C(stage3_c55_s_fa2), .So(stage4_c55_s_fa2), .Co(stage4_c55_c_fa2));
    FA fa_2128(.A(stage3_c55_s_fa3), .B(stage3_c55_s_fa4), .C(stage3_c55_s_fa5), .So(stage4_c55_s_fa3), .Co(stage4_c55_c_fa3));
    FA fa_2129(.A(stage3_c55_c_fa0), .B(stage3_c55_c_fa1), .C(stage3_c55_c_fa2), .So(stage4_c56_s_fa0), .Co(stage4_c56_c_fa0));
    FA fa_2130(.A(stage3_c55_c_fa3), .B(stage3_c55_c_fa4), .C(stage3_c55_c_fa5), .So(stage4_c56_s_fa1), .Co(stage4_c56_c_fa1));
    FA fa_2131(.A(stage3_c56_s_fa0), .B(stage3_c56_s_fa1), .C(stage3_c56_s_fa2), .So(stage4_c56_s_fa2), .Co(stage4_c56_c_fa2));
    FA fa_2132(.A(stage3_c56_s_fa3), .B(stage3_c56_s_fa4), .C(stage3_c56_s_fa5), .So(stage4_c56_s_fa3), .Co(stage4_c56_c_fa3));
    FA fa_2133(.A(stage3_c56_c_fa0), .B(stage3_c56_c_fa1), .C(stage3_c56_c_fa2), .So(stage4_c57_s_fa0), .Co(stage4_c57_c_fa0));
    FA fa_2134(.A(stage3_c56_c_fa3), .B(stage3_c56_c_fa4), .C(stage3_c56_c_fa5), .So(stage4_c57_s_fa1), .Co(stage4_c57_c_fa1));
    FA fa_2135(.A(stage3_c57_s_fa0), .B(stage3_c57_s_fa1), .C(stage3_c57_s_fa2), .So(stage4_c57_s_fa2), .Co(stage4_c57_c_fa2));
    FA fa_2136(.A(stage3_c57_s_fa3), .B(stage3_c57_s_fa4), .C(stage3_c57_s_fa5), .So(stage4_c57_s_fa3), .Co(stage4_c57_c_fa3));
    FA fa_2137(.A(stage3_c57_c_fa0), .B(stage3_c57_c_fa1), .C(stage3_c57_c_fa2), .So(stage4_c58_s_fa0), .Co(stage4_c58_c_fa0));
    FA fa_2138(.A(stage3_c57_c_fa3), .B(stage3_c57_c_fa4), .C(stage3_c57_c_fa5), .So(stage4_c58_s_fa1), .Co(stage4_c58_c_fa1));
    FA fa_2139(.A(stage3_c58_s_fa0), .B(stage3_c58_s_fa1), .C(stage3_c58_s_fa2), .So(stage4_c58_s_fa2), .Co(stage4_c58_c_fa2));
    FA fa_2140(.A(stage3_c58_s_fa3), .B(stage3_c58_s_fa4), .C(stage3_c58_s_fa5), .So(stage4_c58_s_fa3), .Co(stage4_c58_c_fa3));
    FA fa_2141(.A(stage3_c58_c_fa0), .B(stage3_c58_c_fa1), .C(stage3_c58_c_fa2), .So(stage4_c59_s_fa0), .Co(stage4_c59_c_fa0));
    FA fa_2142(.A(stage3_c58_c_fa3), .B(stage3_c58_c_fa4), .C(stage3_c58_c_fa5), .So(stage4_c59_s_fa1), .Co(stage4_c59_c_fa1));
    FA fa_2143(.A(stage3_c59_s_fa0), .B(stage3_c59_s_fa1), .C(stage3_c59_s_fa2), .So(stage4_c59_s_fa2), .Co(stage4_c59_c_fa2));
    FA fa_2144(.A(stage3_c59_s_fa3), .B(stage3_c59_s_fa4), .C(stage3_c59_s_fa5), .So(stage4_c59_s_fa3), .Co(stage4_c59_c_fa3));
    FA fa_2145(.A(stage3_c59_c_fa0), .B(stage3_c59_c_fa1), .C(stage3_c59_c_fa2), .So(stage4_c60_s_fa0), .Co(stage4_c60_c_fa0));
    FA fa_2146(.A(stage3_c59_c_fa3), .B(stage3_c59_c_fa4), .C(stage3_c59_c_fa5), .So(stage4_c60_s_fa1), .Co(stage4_c60_c_fa1));
    FA fa_2147(.A(stage3_c60_s_fa0), .B(stage3_c60_s_fa1), .C(stage3_c60_s_fa2), .So(stage4_c60_s_fa2), .Co(stage4_c60_c_fa2));
    FA fa_2148(.A(stage3_c60_s_fa3), .B(stage3_c60_s_fa4), .C(stage3_c60_s_fa5), .So(stage4_c60_s_fa3), .Co(stage4_c60_c_fa3));
    FA fa_2149(.A(stage3_c60_c_fa0), .B(stage3_c60_c_fa1), .C(stage3_c60_c_fa2), .So(stage4_c61_s_fa0), .Co(stage4_c61_c_fa0));
    FA fa_2150(.A(stage3_c60_c_fa3), .B(stage3_c60_c_fa4), .C(stage3_c60_c_fa5), .So(stage4_c61_s_fa1), .Co(stage4_c61_c_fa1));
    FA fa_2151(.A(stage3_c61_s_fa0), .B(stage3_c61_s_fa1), .C(stage3_c61_s_fa2), .So(stage4_c61_s_fa2), .Co(stage4_c61_c_fa2));
    FA fa_2152(.A(stage3_c61_s_fa3), .B(stage3_c61_s_fa4), .C(stage3_c61_s_fa5), .So(stage4_c61_s_fa3), .Co(stage4_c61_c_fa3));
    FA fa_2153(.A(stage3_c61_c_fa0), .B(stage3_c61_c_fa1), .C(stage3_c61_c_fa2), .So(stage4_c62_s_fa0), .Co(stage4_c62_c_fa0));
    FA fa_2154(.A(stage3_c61_c_fa3), .B(stage3_c61_c_fa4), .C(stage3_c61_c_fa5), .So(stage4_c62_s_fa1), .Co(stage4_c62_c_fa1));
    FA fa_2155(.A(stage3_c62_s_fa0), .B(stage3_c62_s_fa1), .C(stage3_c62_s_fa2), .So(stage4_c62_s_fa2), .Co(stage4_c62_c_fa2));
    FA fa_2156(.A(stage3_c62_s_fa3), .B(stage3_c62_s_fa4), .C(stage3_c62_s_fa5), .So(stage4_c62_s_fa3), .Co(stage4_c62_c_fa3));
    FA fa_2157(.A(stage3_c62_c_fa0), .B(stage3_c62_c_fa1), .C(stage3_c62_c_fa2), .So(stage4_c63_s_fa0), .Co(stage4_c63_c_fa0));
    FA fa_2158(.A(stage3_c62_c_fa3), .B(stage3_c62_c_fa4), .C(stage3_c62_c_fa5), .So(stage4_c63_s_fa1), .Co(stage4_c63_c_fa1));
    FA fa_2159(.A(stage3_c63_s_fa0), .B(stage3_c63_s_fa1), .C(stage3_c63_s_fa2), .So(stage4_c63_s_fa2), .Co(stage4_c63_c_fa2));
    FA fa_2160(.A(stage3_c63_s_fa3), .B(stage3_c63_s_fa4), .C(stage3_c63_s_fa5), .So(stage4_c63_s_fa3), .Co(stage4_c63_c_fa3));
    FA fa_2161(.A(stage3_c63_c_fa0), .B(stage3_c63_c_fa1), .C(stage3_c63_c_fa2), .So(stage4_c64_s_fa0), .Co(stage4_c64_c_fa0));
    FA fa_2162(.A(stage3_c63_c_fa3), .B(stage3_c63_c_fa4), .C(stage3_c63_c_fa5), .So(stage4_c64_s_fa1), .Co(stage4_c64_c_fa1));
    FA fa_2163(.A(stage3_c64_s_fa0), .B(stage3_c64_s_fa1), .C(stage3_c64_s_fa2), .So(stage4_c64_s_fa2), .Co(stage4_c64_c_fa2));
    FA fa_2164(.A(stage3_c64_s_fa3), .B(stage3_c64_s_fa4), .C(stage3_c64_s_fa5), .So(stage4_c64_s_fa3), .Co(stage4_c64_c_fa3));
    FA fa_2165(.A(stage3_c64_c_fa0), .B(stage3_c64_c_fa1), .C(stage3_c64_c_fa2), .So(stage4_c65_s_fa0), .Co(stage4_c65_c_fa0));
    FA fa_2166(.A(stage3_c64_c_fa3), .B(stage3_c64_c_fa4), .C(stage3_c64_c_fa5), .So(stage4_c65_s_fa1), .Co(stage4_c65_c_fa1));
    FA fa_2167(.A(stage3_c65_s_fa0), .B(stage3_c65_s_fa1), .C(stage3_c65_s_fa2), .So(stage4_c65_s_fa2), .Co(stage4_c65_c_fa2));
    FA fa_2168(.A(stage3_c65_s_fa3), .B(stage3_c65_s_fa4), .C(stage3_c65_s_fa5), .So(stage4_c65_s_fa3), .Co(stage4_c65_c_fa3));
    FA fa_2169(.A(stage3_c65_c_fa0), .B(stage3_c65_c_fa1), .C(stage3_c65_c_fa2), .So(stage4_c66_s_fa0), .Co(stage4_c66_c_fa0));
    FA fa_2170(.A(stage3_c65_c_fa3), .B(stage3_c65_c_fa4), .C(stage3_c65_c_fa5), .So(stage4_c66_s_fa1), .Co(stage4_c66_c_fa1));
    FA fa_2171(.A(stage3_c66_s_fa0), .B(stage3_c66_s_fa1), .C(stage3_c66_s_fa2), .So(stage4_c66_s_fa2), .Co(stage4_c66_c_fa2));
    FA fa_2172(.A(stage3_c66_s_fa3), .B(stage3_c66_s_fa4), .C(stage3_c66_s_fa5), .So(stage4_c66_s_fa3), .Co(stage4_c66_c_fa3));
    FA fa_2173(.A(stage3_c66_c_fa0), .B(stage3_c66_c_fa1), .C(stage3_c66_c_fa2), .So(stage4_c67_s_fa0), .Co(stage4_c67_c_fa0));
    FA fa_2174(.A(stage3_c66_c_fa3), .B(stage3_c66_c_fa4), .C(stage3_c66_c_fa5), .So(stage4_c67_s_fa1), .Co(stage4_c67_c_fa1));
    FA fa_2175(.A(stage3_c67_s_fa0), .B(stage3_c67_s_fa1), .C(stage3_c67_s_fa2), .So(stage4_c67_s_fa2), .Co(stage4_c67_c_fa2));
    FA fa_2176(.A(stage3_c67_s_fa3), .B(stage3_c67_s_fa4), .C(stage3_c67_s_fa5), .So(stage4_c67_s_fa3), .Co(stage4_c67_c_fa3));
    FA fa_2177(.A(stage3_c67_c_fa0), .B(stage3_c67_c_fa1), .C(stage3_c67_c_fa2), .So(stage4_c68_s_fa0), .Co(stage4_c68_c_fa0));
    FA fa_2178(.A(stage3_c67_c_fa3), .B(stage3_c67_c_fa4), .C(stage3_c67_c_fa5), .So(stage4_c68_s_fa1), .Co(stage4_c68_c_fa1));
    FA fa_2179(.A(stage3_c68_s_fa0), .B(stage3_c68_s_fa1), .C(stage3_c68_s_fa2), .So(stage4_c68_s_fa2), .Co(stage4_c68_c_fa2));
    FA fa_2180(.A(stage3_c68_s_fa3), .B(stage3_c68_s_fa4), .C(stage3_c68_s_fa5), .So(stage4_c68_s_fa3), .Co(stage4_c68_c_fa3));
    FA fa_2181(.A(stage3_c68_c_fa0), .B(stage3_c68_c_fa1), .C(stage3_c68_c_fa2), .So(stage4_c69_s_fa0), .Co(stage4_c69_c_fa0));
    FA fa_2182(.A(stage3_c68_c_fa3), .B(stage3_c68_c_fa4), .C(stage3_c68_c_fa5), .So(stage4_c69_s_fa1), .Co(stage4_c69_c_fa1));
    FA fa_2183(.A(stage3_c69_s_fa0), .B(stage3_c69_s_fa1), .C(stage3_c69_s_fa2), .So(stage4_c69_s_fa2), .Co(stage4_c69_c_fa2));
    FA fa_2184(.A(stage3_c69_s_fa3), .B(stage3_c69_s_fa4), .C(stage3_c69_s_fa5), .So(stage4_c69_s_fa3), .Co(stage4_c69_c_fa3));
    FA fa_2185(.A(stage3_c69_c_fa0), .B(stage3_c69_c_fa1), .C(stage3_c69_c_fa2), .So(stage4_c70_s_fa0), .Co(stage4_c70_c_fa0));
    FA fa_2186(.A(stage3_c69_c_fa3), .B(stage3_c69_c_fa4), .C(stage3_c69_c_fa5), .So(stage4_c70_s_fa1), .Co(stage4_c70_c_fa1));
    FA fa_2187(.A(stage3_c70_s_fa0), .B(stage3_c70_s_fa1), .C(stage3_c70_s_fa2), .So(stage4_c70_s_fa2), .Co(stage4_c70_c_fa2));
    FA fa_2188(.A(stage3_c70_s_fa3), .B(stage3_c70_s_fa4), .C(stage3_c70_s_fa5), .So(stage4_c70_s_fa3), .Co(stage4_c70_c_fa3));
    FA fa_2189(.A(stage3_c70_c_fa0), .B(stage3_c70_c_fa1), .C(stage3_c70_c_fa2), .So(stage4_c71_s_fa0), .Co(stage4_c71_c_fa0));
    FA fa_2190(.A(stage3_c70_c_fa3), .B(stage3_c70_c_fa4), .C(stage3_c70_c_fa5), .So(stage4_c71_s_fa1), .Co(stage4_c71_c_fa1));
    FA fa_2191(.A(stage3_c71_s_fa0), .B(stage3_c71_s_fa1), .C(stage3_c71_s_fa2), .So(stage4_c71_s_fa2), .Co(stage4_c71_c_fa2));
    FA fa_2192(.A(stage3_c71_s_fa3), .B(stage3_c71_s_fa4), .C(stage3_c71_s_fa5), .So(stage4_c71_s_fa3), .Co(stage4_c71_c_fa3));
    FA fa_2193(.A(stage3_c71_c_fa0), .B(stage3_c71_c_fa1), .C(stage3_c71_c_fa2), .So(stage4_c72_s_fa0), .Co(stage4_c72_c_fa0));
    FA fa_2194(.A(stage3_c71_c_fa3), .B(stage3_c71_c_fa4), .C(stage3_c71_c_fa5), .So(stage4_c72_s_fa1), .Co(stage4_c72_c_fa1));
    FA fa_2195(.A(stage3_c72_s_fa0), .B(stage3_c72_s_fa1), .C(stage3_c72_s_fa2), .So(stage4_c72_s_fa2), .Co(stage4_c72_c_fa2));
    FA fa_2196(.A(stage3_c72_s_fa3), .B(stage3_c72_s_fa4), .C(stage3_c72_s_fa5), .So(stage4_c72_s_fa3), .Co(stage4_c72_c_fa3));
    FA fa_2197(.A(stage3_c72_c_fa0), .B(stage3_c72_c_fa1), .C(stage3_c72_c_fa2), .So(stage4_c73_s_fa0), .Co(stage4_c73_c_fa0));
    FA fa_2198(.A(stage3_c72_c_fa3), .B(stage3_c72_c_fa4), .C(stage3_c72_c_fa5), .So(stage4_c73_s_fa1), .Co(stage4_c73_c_fa1));
    FA fa_2199(.A(stage3_c73_s_fa0), .B(stage3_c73_s_fa1), .C(stage3_c73_s_fa2), .So(stage4_c73_s_fa2), .Co(stage4_c73_c_fa2));
    FA fa_2200(.A(stage3_c73_s_fa3), .B(stage3_c73_s_fa4), .C(stage3_c73_s_fa5), .So(stage4_c73_s_fa3), .Co(stage4_c73_c_fa3));
    FA fa_2201(.A(stage3_c73_c_fa0), .B(stage3_c73_c_fa1), .C(stage3_c73_c_fa2), .So(stage4_c74_s_fa0), .Co(stage4_c74_c_fa0));
    FA fa_2202(.A(stage3_c73_c_fa3), .B(stage3_c73_c_fa4), .C(stage3_c73_c_fa5), .So(stage4_c74_s_fa1), .Co(stage4_c74_c_fa1));
    FA fa_2203(.A(stage3_c74_s_fa0), .B(stage3_c74_s_fa1), .C(stage3_c74_s_fa2), .So(stage4_c74_s_fa2), .Co(stage4_c74_c_fa2));
    FA fa_2204(.A(stage3_c74_s_fa3), .B(stage3_c74_s_fa4), .C(stage3_c74_s_fa5), .So(stage4_c74_s_fa3), .Co(stage4_c74_c_fa3));
    FA fa_2205(.A(stage3_c74_c_fa0), .B(stage3_c74_c_fa1), .C(stage3_c74_c_fa2), .So(stage4_c75_s_fa0), .Co(stage4_c75_c_fa0));
    FA fa_2206(.A(stage3_c74_c_fa3), .B(stage3_c74_c_fa4), .C(stage3_c74_c_fa5), .So(stage4_c75_s_fa1), .Co(stage4_c75_c_fa1));
    FA fa_2207(.A(stage3_c75_s_fa0), .B(stage3_c75_s_fa1), .C(stage3_c75_s_fa2), .So(stage4_c75_s_fa2), .Co(stage4_c75_c_fa2));
    FA fa_2208(.A(stage3_c75_s_fa3), .B(stage3_c75_s_fa4), .C(stage3_c75_s_fa5), .So(stage4_c75_s_fa3), .Co(stage4_c75_c_fa3));
    FA fa_2209(.A(stage3_c75_c_fa0), .B(stage3_c75_c_fa1), .C(stage3_c75_c_fa2), .So(stage4_c76_s_fa0), .Co(stage4_c76_c_fa0));
    FA fa_2210(.A(stage3_c75_c_fa3), .B(stage3_c75_c_fa4), .C(stage3_c75_c_fa5), .So(stage4_c76_s_fa1), .Co(stage4_c76_c_fa1));
    FA fa_2211(.A(stage3_c76_s_fa0), .B(stage3_c76_s_fa1), .C(stage3_c76_s_fa2), .So(stage4_c76_s_fa2), .Co(stage4_c76_c_fa2));
    FA fa_2212(.A(stage3_c76_s_fa3), .B(stage3_c76_s_fa4), .C(stage3_c76_s_ha0), .So(stage4_c76_s_fa3), .Co(stage4_c76_c_fa3));
    FA fa_2213(.A(stage3_c76_c_fa0), .B(stage3_c76_c_fa1), .C(stage3_c76_c_fa2), .So(stage4_c77_s_fa0), .Co(stage4_c77_c_fa0));
    FA fa_2214(.A(stage3_c76_c_fa3), .B(stage3_c76_c_fa4), .C(stage3_c76_c_ha0), .So(stage4_c77_s_fa1), .Co(stage4_c77_c_fa1));
    FA fa_2215(.A(stage3_c77_s_fa0), .B(stage3_c77_s_fa1), .C(stage3_c77_s_fa2), .So(stage4_c77_s_fa2), .Co(stage4_c77_c_fa2));
    FA fa_2216(.A(stage3_c77_s_fa3), .B(stage3_c77_s_fa4), .C(stage2_c77_s_fa7), .So(stage4_c77_s_fa3), .Co(stage4_c77_c_fa3));
    FA fa_2217(.A(stage3_c77_c_fa0), .B(stage3_c77_c_fa1), .C(stage3_c77_c_fa2), .So(stage4_c78_s_fa0), .Co(stage4_c78_c_fa0));
    FA fa_2218(.A(stage3_c77_c_fa3), .B(stage3_c77_c_fa4), .C(stage3_c78_s_fa0), .So(stage4_c78_s_fa1), .Co(stage4_c78_c_fa1));
    FA fa_2219(.A(stage3_c78_s_fa1), .B(stage3_c78_s_fa2), .C(stage3_c78_s_fa3), .So(stage4_c78_s_fa2), .Co(stage4_c78_c_fa2));
    HA ha_125(.A(stage3_c78_s_fa4), .B(stage2_c78_s_fa7), .So(stage4_c78_s_ha0), .Co(stage4_c78_c_ha0));
    FA fa_2220(.A(stage3_c78_c_fa0), .B(stage3_c78_c_fa1), .C(stage3_c78_c_fa2), .So(stage4_c79_s_fa0), .Co(stage4_c79_c_fa0));
    FA fa_2221(.A(stage3_c78_c_fa3), .B(stage3_c78_c_fa4), .C(stage3_c79_s_fa0), .So(stage4_c79_s_fa1), .Co(stage4_c79_c_fa1));
    FA fa_2222(.A(stage3_c79_s_fa1), .B(stage3_c79_s_fa2), .C(stage3_c79_s_fa3), .So(stage4_c79_s_fa2), .Co(stage4_c79_c_fa2));
    HA ha_126(.A(stage3_c79_s_fa4), .B(stage1_c79_s_fa10), .So(stage4_c79_s_ha0), .Co(stage4_c79_c_ha0));
    FA fa_2223(.A(stage3_c79_c_fa0), .B(stage3_c79_c_fa1), .C(stage3_c79_c_fa2), .So(stage4_c80_s_fa0), .Co(stage4_c80_c_fa0));
    FA fa_2224(.A(stage3_c79_c_fa3), .B(stage3_c79_c_fa4), .C(stage3_c80_s_fa0), .So(stage4_c80_s_fa1), .Co(stage4_c80_c_fa1));
    FA fa_2225(.A(stage3_c80_s_fa1), .B(stage3_c80_s_fa2), .C(stage3_c80_s_fa3), .So(stage4_c80_s_fa2), .Co(stage4_c80_c_fa2));
    FA fa_2226(.A(stage3_c80_c_fa0), .B(stage3_c80_c_fa1), .C(stage3_c80_c_fa2), .So(stage4_c81_s_fa0), .Co(stage4_c81_c_fa0));
    FA fa_2227(.A(stage3_c80_c_fa3), .B(stage3_c80_c_fa4), .C(stage3_c81_s_fa0), .So(stage4_c81_s_fa1), .Co(stage4_c81_c_fa1));
    FA fa_2228(.A(stage3_c81_s_fa1), .B(stage3_c81_s_fa2), .C(stage3_c81_s_fa3), .So(stage4_c81_s_fa2), .Co(stage4_c81_c_fa2));
    FA fa_2229(.A(stage3_c81_c_fa0), .B(stage3_c81_c_fa1), .C(stage3_c81_c_fa2), .So(stage4_c82_s_fa0), .Co(stage4_c82_c_fa0));
    FA fa_2230(.A(stage3_c81_c_fa3), .B(stage3_c81_c_fa4), .C(stage3_c82_s_fa0), .So(stage4_c82_s_fa1), .Co(stage4_c82_c_fa1));
    FA fa_2231(.A(stage3_c82_s_fa1), .B(stage3_c82_s_fa2), .C(stage3_c82_s_fa3), .So(stage4_c82_s_fa2), .Co(stage4_c82_c_fa2));
    FA fa_2232(.A(stage3_c82_c_fa0), .B(stage3_c82_c_fa1), .C(stage3_c82_c_fa2), .So(stage4_c83_s_fa0), .Co(stage4_c83_c_fa0));
    FA fa_2233(.A(stage3_c82_c_fa3), .B(stage3_c82_c_ha0), .C(stage3_c83_s_fa0), .So(stage4_c83_s_fa1), .Co(stage4_c83_c_fa1));
    FA fa_2234(.A(stage3_c83_s_fa1), .B(stage3_c83_s_fa2), .C(stage3_c83_s_fa3), .So(stage4_c83_s_fa2), .Co(stage4_c83_c_fa2));
    FA fa_2235(.A(stage3_c83_c_fa0), .B(stage3_c83_c_fa1), .C(stage3_c83_c_fa2), .So(stage4_c84_s_fa0), .Co(stage4_c84_c_fa0));
    FA fa_2236(.A(stage3_c83_c_fa3), .B(stage3_c83_c_ha0), .C(stage3_c84_s_fa0), .So(stage4_c84_s_fa1), .Co(stage4_c84_c_fa1));
    FA fa_2237(.A(stage3_c84_s_fa1), .B(stage3_c84_s_fa2), .C(stage3_c84_s_fa3), .So(stage4_c84_s_fa2), .Co(stage4_c84_c_fa2));
    FA fa_2238(.A(stage3_c84_c_fa0), .B(stage3_c84_c_fa1), .C(stage3_c84_c_fa2), .So(stage4_c85_s_fa0), .Co(stage4_c85_c_fa0));
    FA fa_2239(.A(stage3_c84_c_fa3), .B(stage3_c84_c_ha0), .C(stage3_c85_s_fa0), .So(stage4_c85_s_fa1), .Co(stage4_c85_c_fa1));
    FA fa_2240(.A(stage3_c85_s_fa1), .B(stage3_c85_s_fa2), .C(stage3_c85_s_fa3), .So(stage4_c85_s_fa2), .Co(stage4_c85_c_fa2));
    FA fa_2241(.A(stage3_c85_c_fa0), .B(stage3_c85_c_fa1), .C(stage3_c85_c_fa2), .So(stage4_c86_s_fa0), .Co(stage4_c86_c_fa0));
    FA fa_2242(.A(stage3_c85_c_fa3), .B(stage3_c86_s_fa0), .C(stage3_c86_s_fa1), .So(stage4_c86_s_fa1), .Co(stage4_c86_c_fa1));
    HA ha_127(.A(stage3_c86_s_fa2), .B(stage3_c86_s_fa3), .So(stage4_c86_s_ha0), .Co(stage4_c86_c_ha0));
    FA fa_2243(.A(stage3_c86_c_fa0), .B(stage3_c86_c_fa1), .C(stage3_c86_c_fa2), .So(stage4_c87_s_fa0), .Co(stage4_c87_c_fa0));
    FA fa_2244(.A(stage3_c86_c_fa3), .B(stage3_c87_s_fa0), .C(stage3_c87_s_fa1), .So(stage4_c87_s_fa1), .Co(stage4_c87_c_fa1));
    HA ha_128(.A(stage3_c87_s_fa2), .B(stage3_c87_s_fa3), .So(stage4_c87_s_ha0), .Co(stage4_c87_c_ha0));
    FA fa_2245(.A(stage3_c87_c_fa0), .B(stage3_c87_c_fa1), .C(stage3_c87_c_fa2), .So(stage4_c88_s_fa0), .Co(stage4_c88_c_fa0));
    FA fa_2246(.A(stage3_c87_c_fa3), .B(stage3_c88_s_fa0), .C(stage3_c88_s_fa1), .So(stage4_c88_s_fa1), .Co(stage4_c88_c_fa1));
    HA ha_129(.A(stage3_c88_s_fa2), .B(stage3_c88_s_fa3), .So(stage4_c88_s_ha0), .Co(stage4_c88_c_ha0));
    FA fa_2247(.A(stage3_c88_c_fa0), .B(stage3_c88_c_fa1), .C(stage3_c88_c_fa2), .So(stage4_c89_s_fa0), .Co(stage4_c89_c_fa0));
    FA fa_2248(.A(stage3_c88_c_fa3), .B(stage3_c89_s_fa0), .C(stage3_c89_s_fa1), .So(stage4_c89_s_fa1), .Co(stage4_c89_c_fa1));
    HA ha_130(.A(stage3_c89_s_fa2), .B(stage3_c89_s_ha0), .So(stage4_c89_s_ha0), .Co(stage4_c89_c_ha0));
    FA fa_2249(.A(stage3_c89_c_fa0), .B(stage3_c89_c_fa1), .C(stage3_c89_c_fa2), .So(stage4_c90_s_fa0), .Co(stage4_c90_c_fa0));
    FA fa_2250(.A(stage3_c89_c_ha0), .B(stage3_c90_s_fa0), .C(stage3_c90_s_fa1), .So(stage4_c90_s_fa1), .Co(stage4_c90_c_fa1));
    HA ha_131(.A(stage3_c90_s_fa2), .B(stage3_c90_s_ha0), .So(stage4_c90_s_ha0), .Co(stage4_c90_c_ha0));
    FA fa_2251(.A(stage3_c90_c_fa0), .B(stage3_c90_c_fa1), .C(stage3_c90_c_fa2), .So(stage4_c91_s_fa0), .Co(stage4_c91_c_fa0));
    FA fa_2252(.A(stage3_c90_c_ha0), .B(stage3_c91_s_fa0), .C(stage3_c91_s_fa1), .So(stage4_c91_s_fa1), .Co(stage4_c91_c_fa1));
    HA ha_132(.A(stage3_c91_s_fa2), .B(stage2_c91_s_ha0), .So(stage4_c91_s_ha0), .Co(stage4_c91_c_ha0));
    FA fa_2253(.A(stage3_c91_c_fa0), .B(stage3_c91_c_fa1), .C(stage3_c91_c_fa2), .So(stage4_c92_s_fa0), .Co(stage4_c92_c_fa0));
    FA fa_2254(.A(stage3_c92_s_fa0), .B(stage3_c92_s_fa1), .C(stage3_c92_s_fa2), .So(stage4_c92_s_fa1), .Co(stage4_c92_c_fa1));
    FA fa_2255(.A(stage3_c92_c_fa0), .B(stage3_c92_c_fa1), .C(stage3_c92_c_fa2), .So(stage4_c93_s_fa0), .Co(stage4_c93_c_fa0));
    FA fa_2256(.A(stage3_c93_s_fa0), .B(stage3_c93_s_fa1), .C(stage3_c93_s_fa2), .So(stage4_c93_s_fa1), .Co(stage4_c93_c_fa1));
    FA fa_2257(.A(stage3_c93_c_fa0), .B(stage3_c93_c_fa1), .C(stage3_c93_c_fa2), .So(stage4_c94_s_fa0), .Co(stage4_c94_c_fa0));
    FA fa_2258(.A(stage3_c94_s_fa0), .B(stage3_c94_s_fa1), .C(stage3_c94_s_fa2), .So(stage4_c94_s_fa1), .Co(stage4_c94_c_fa1));
    FA fa_2259(.A(stage3_c94_c_fa0), .B(stage3_c94_c_fa1), .C(stage3_c94_c_fa2), .So(stage4_c95_s_fa0), .Co(stage4_c95_c_fa0));
    FA fa_2260(.A(stage3_c95_s_fa0), .B(stage3_c95_s_fa1), .C(stage3_c95_s_ha0), .So(stage4_c95_s_fa1), .Co(stage4_c95_c_fa1));
    FA fa_2261(.A(stage3_c95_c_fa0), .B(stage3_c95_c_fa1), .C(stage3_c95_c_ha0), .So(stage4_c96_s_fa0), .Co(stage4_c96_c_fa0));
    FA fa_2262(.A(stage3_c96_s_fa0), .B(stage3_c96_s_fa1), .C(stage3_c96_s_ha0), .So(stage4_c96_s_fa1), .Co(stage4_c96_c_fa1));
    FA fa_2263(.A(stage3_c96_c_fa0), .B(stage3_c96_c_fa1), .C(stage3_c96_c_ha0), .So(stage4_c97_s_fa0), .Co(stage4_c97_c_fa0));
    FA fa_2264(.A(stage3_c97_s_fa0), .B(stage3_c97_s_fa1), .C(stage3_c97_s_ha0), .So(stage4_c97_s_fa1), .Co(stage4_c97_c_fa1));
    FA fa_2265(.A(stage3_c97_c_fa0), .B(stage3_c97_c_fa1), .C(stage3_c97_c_ha0), .So(stage4_c98_s_fa0), .Co(stage4_c98_c_fa0));
    FA fa_2266(.A(stage3_c98_s_fa0), .B(stage3_c98_s_fa1), .C(stage1_c98_s_ha0), .So(stage4_c98_s_fa1), .Co(stage4_c98_c_fa1));
    FA fa_2267(.A(stage3_c98_c_fa0), .B(stage3_c98_c_fa1), .C(stage3_c99_s_fa0), .So(stage4_c99_s_fa0), .Co(stage4_c99_c_fa0));
    HA ha_133(.A(stage3_c99_s_fa1), .B(stage0_r71_c28), .So(stage4_c99_s_ha0), .Co(stage4_c99_c_ha0));
    FA fa_2268(.A(stage3_c99_c_fa0), .B(stage3_c99_c_fa1), .C(stage3_c100_s_fa0), .So(stage4_c100_s_fa0), .Co(stage4_c100_c_fa0));
    FA fa_2269(.A(stage3_c100_c_fa0), .B(stage3_c100_c_fa1), .C(stage3_c101_s_fa0), .So(stage4_c101_s_fa0), .Co(stage4_c101_c_fa0));
    FA fa_2270(.A(stage3_c101_c_fa0), .B(stage3_c101_c_fa1), .C(stage3_c102_s_fa0), .So(stage4_c102_s_fa0), .Co(stage4_c102_c_fa0));
    FA fa_2271(.A(stage3_c102_c_fa0), .B(stage3_c102_c_fa1), .C(stage3_c103_s_fa0), .So(stage4_c103_s_fa0), .Co(stage4_c103_c_fa0));
    FA fa_2272(.A(stage3_c103_c_fa0), .B(stage3_c103_c_ha0), .C(stage3_c104_s_fa0), .So(stage4_c104_s_fa0), .Co(stage4_c104_c_fa0));
    FA fa_2273(.A(stage3_c104_c_fa0), .B(stage3_c105_s_fa0), .C(stage2_c105_s_fa1), .So(stage4_c105_s_fa0), .Co(stage4_c105_c_fa0));
    FA fa_2274(.A(stage3_c105_c_fa0), .B(stage3_c106_s_fa0), .C(stage1_c106_s_fa1), .So(stage4_c106_s_fa0), .Co(stage4_c106_c_fa0));
    HA ha_134(.A(stage3_c106_c_fa0), .B(stage3_c107_s_fa0), .So(stage4_c107_s_ha0), .Co(stage4_c107_c_ha0));
    HA ha_135(.A(stage3_c107_c_fa0), .B(stage3_c108_s_fa0), .So(stage4_c108_s_ha0), .Co(stage4_c108_c_ha0));
    HA ha_136(.A(stage3_c108_c_fa0), .B(stage3_c109_s_ha0), .So(stage4_c109_s_ha0), .Co(stage4_c109_c_ha0));
    HA ha_137(.A(stage3_c109_c_ha0), .B(stage3_c110_s_ha0), .So(stage4_c110_s_ha0), .Co(stage4_c110_c_ha0));
    HA ha_138(.A(stage3_c110_c_ha0), .B(stage3_c111_s_ha0), .So(stage4_c111_s_ha0), .Co(stage4_c111_c_ha0));
    HA ha_139(.A(stage3_c111_c_ha0), .B(stage2_c111_c_ha0), .So(stage4_c112_s_ha0), .Co(stage4_c112_c_ha0));
    HA ha_140(.A(stage4_c4_c_ha0), .B(stage4_c5_s_ha0), .So(stage5_c5_s_ha0), .Co(stage5_c5_c_ha0));
    HA ha_141(.A(stage4_c5_c_ha0), .B(stage4_c6_s_ha0), .So(stage5_c6_s_ha0), .Co(stage5_c6_c_ha0));
    HA ha_142(.A(stage4_c6_c_ha0), .B(stage4_c7_s_fa0), .So(stage5_c7_s_ha0), .Co(stage5_c7_c_ha0));
    HA ha_143(.A(stage4_c7_c_fa0), .B(stage4_c8_s_fa0), .So(stage5_c8_s_ha0), .Co(stage5_c8_c_ha0));
    HA ha_144(.A(stage4_c8_c_fa0), .B(stage4_c9_s_fa0), .So(stage5_c9_s_ha0), .Co(stage5_c9_c_ha0));
    FA fa_2275(.A(stage4_c9_c_fa0), .B(stage4_c10_s_fa0), .C(stage3_c10_s_ha0), .So(stage5_c10_s_fa0), .Co(stage5_c10_c_fa0));
    FA fa_2276(.A(stage4_c10_c_fa0), .B(stage4_c11_s_fa0), .C(stage3_c11_s_ha0), .So(stage5_c11_s_fa0), .Co(stage5_c11_c_fa0));
    FA fa_2277(.A(stage4_c11_c_fa0), .B(stage4_c12_s_fa0), .C(stage3_c12_s_fa1), .So(stage5_c12_s_fa0), .Co(stage5_c12_c_fa0));
    FA fa_2278(.A(stage4_c12_c_fa0), .B(stage4_c13_s_fa0), .C(stage3_c13_s_fa1), .So(stage5_c13_s_fa0), .Co(stage5_c13_c_fa0));
    FA fa_2279(.A(stage4_c13_c_fa0), .B(stage4_c14_s_fa0), .C(stage4_c14_s_ha0), .So(stage5_c14_s_fa0), .Co(stage5_c14_c_fa0));
    FA fa_2280(.A(stage4_c14_c_fa0), .B(stage4_c14_c_ha0), .C(stage4_c15_s_fa0), .So(stage5_c15_s_fa0), .Co(stage5_c15_c_fa0));
    FA fa_2281(.A(stage4_c15_c_fa0), .B(stage4_c15_c_ha0), .C(stage4_c16_s_fa0), .So(stage5_c16_s_fa0), .Co(stage5_c16_c_fa0));
    FA fa_2282(.A(stage4_c16_c_fa0), .B(stage4_c16_c_ha0), .C(stage4_c17_s_fa0), .So(stage5_c17_s_fa0), .Co(stage5_c17_c_fa0));
    FA fa_2283(.A(stage4_c17_c_fa0), .B(stage4_c17_c_fa1), .C(stage4_c18_s_fa0), .So(stage5_c18_s_fa0), .Co(stage5_c18_c_fa0));
    FA fa_2284(.A(stage4_c18_c_fa0), .B(stage4_c18_c_fa1), .C(stage4_c19_s_fa0), .So(stage5_c19_s_fa0), .Co(stage5_c19_c_fa0));
    FA fa_2285(.A(stage4_c19_c_fa0), .B(stage4_c19_c_fa1), .C(stage4_c20_s_fa0), .So(stage5_c20_s_fa0), .Co(stage5_c20_c_fa0));
    FA fa_2286(.A(stage4_c20_c_fa0), .B(stage4_c20_c_fa1), .C(stage4_c21_s_fa0), .So(stage5_c21_s_fa0), .Co(stage5_c21_c_fa0));
    HA ha_145(.A(stage4_c21_s_fa1), .B(stage2_c21_s_fa4), .So(stage5_c21_s_ha0), .Co(stage5_c21_c_ha0));
    FA fa_2287(.A(stage4_c21_c_fa0), .B(stage4_c21_c_fa1), .C(stage4_c22_s_fa0), .So(stage5_c22_s_fa0), .Co(stage5_c22_c_fa0));
    HA ha_146(.A(stage4_c22_s_fa1), .B(stage2_c22_s_fa4), .So(stage5_c22_s_ha0), .Co(stage5_c22_c_ha0));
    FA fa_2288(.A(stage4_c22_c_fa0), .B(stage4_c22_c_fa1), .C(stage4_c23_s_fa0), .So(stage5_c23_s_fa0), .Co(stage5_c23_c_fa0));
    HA ha_147(.A(stage4_c23_s_fa1), .B(stage3_c23_s_ha0), .So(stage5_c23_s_ha0), .Co(stage5_c23_c_ha0));
    FA fa_2289(.A(stage4_c23_c_fa0), .B(stage4_c23_c_fa1), .C(stage4_c24_s_fa0), .So(stage5_c24_s_fa0), .Co(stage5_c24_c_fa0));
    HA ha_148(.A(stage4_c24_s_fa1), .B(stage4_c24_s_ha0), .So(stage5_c24_s_ha0), .Co(stage5_c24_c_ha0));
    FA fa_2290(.A(stage4_c24_c_fa0), .B(stage4_c24_c_fa1), .C(stage4_c24_c_ha0), .So(stage5_c25_s_fa0), .Co(stage5_c25_c_fa0));
    FA fa_2291(.A(stage4_c25_s_fa0), .B(stage4_c25_s_fa1), .C(stage4_c25_s_ha0), .So(stage5_c25_s_fa1), .Co(stage5_c25_c_fa1));
    FA fa_2292(.A(stage4_c25_c_fa0), .B(stage4_c25_c_fa1), .C(stage4_c25_c_ha0), .So(stage5_c26_s_fa0), .Co(stage5_c26_c_fa0));
    FA fa_2293(.A(stage4_c26_s_fa0), .B(stage4_c26_s_fa1), .C(stage4_c26_s_ha0), .So(stage5_c26_s_fa1), .Co(stage5_c26_c_fa1));
    FA fa_2294(.A(stage4_c26_c_fa0), .B(stage4_c26_c_fa1), .C(stage4_c26_c_ha0), .So(stage5_c27_s_fa0), .Co(stage5_c27_c_fa0));
    FA fa_2295(.A(stage4_c27_s_fa0), .B(stage4_c27_s_fa1), .C(stage4_c27_s_fa2), .So(stage5_c27_s_fa1), .Co(stage5_c27_c_fa1));
    FA fa_2296(.A(stage4_c27_c_fa0), .B(stage4_c27_c_fa1), .C(stage4_c27_c_fa2), .So(stage5_c28_s_fa0), .Co(stage5_c28_c_fa0));
    FA fa_2297(.A(stage4_c28_s_fa0), .B(stage4_c28_s_fa1), .C(stage4_c28_s_fa2), .So(stage5_c28_s_fa1), .Co(stage5_c28_c_fa1));
    FA fa_2298(.A(stage4_c28_c_fa0), .B(stage4_c28_c_fa1), .C(stage4_c28_c_fa2), .So(stage5_c29_s_fa0), .Co(stage5_c29_c_fa0));
    FA fa_2299(.A(stage4_c29_s_fa0), .B(stage4_c29_s_fa1), .C(stage4_c29_s_fa2), .So(stage5_c29_s_fa1), .Co(stage5_c29_c_fa1));
    FA fa_2300(.A(stage4_c29_c_fa0), .B(stage4_c29_c_fa1), .C(stage4_c29_c_fa2), .So(stage5_c30_s_fa0), .Co(stage5_c30_c_fa0));
    FA fa_2301(.A(stage4_c30_s_fa0), .B(stage4_c30_s_fa1), .C(stage4_c30_s_fa2), .So(stage5_c30_s_fa1), .Co(stage5_c30_c_fa1));
    FA fa_2302(.A(stage4_c30_c_fa0), .B(stage4_c30_c_fa1), .C(stage4_c30_c_fa2), .So(stage5_c31_s_fa0), .Co(stage5_c31_c_fa0));
    FA fa_2303(.A(stage4_c31_s_fa0), .B(stage4_c31_s_fa1), .C(stage4_c31_s_fa2), .So(stage5_c31_s_fa1), .Co(stage5_c31_c_fa1));
    FA fa_2304(.A(stage4_c31_c_fa0), .B(stage4_c31_c_fa1), .C(stage4_c31_c_fa2), .So(stage5_c32_s_fa0), .Co(stage5_c32_c_fa0));
    FA fa_2305(.A(stage4_c32_s_fa0), .B(stage4_c32_s_fa1), .C(stage4_c32_s_fa2), .So(stage5_c32_s_fa1), .Co(stage5_c32_c_fa1));
    FA fa_2306(.A(stage4_c32_c_fa0), .B(stage4_c32_c_fa1), .C(stage4_c32_c_fa2), .So(stage5_c33_s_fa0), .Co(stage5_c33_c_fa0));
    FA fa_2307(.A(stage4_c33_s_fa0), .B(stage4_c33_s_fa1), .C(stage4_c33_s_fa2), .So(stage5_c33_s_fa1), .Co(stage5_c33_c_fa1));
    FA fa_2308(.A(stage4_c33_c_fa0), .B(stage4_c33_c_fa1), .C(stage4_c33_c_fa2), .So(stage5_c34_s_fa0), .Co(stage5_c34_c_fa0));
    FA fa_2309(.A(stage4_c34_s_fa0), .B(stage4_c34_s_fa1), .C(stage4_c34_s_fa2), .So(stage5_c34_s_fa1), .Co(stage5_c34_c_fa1));
    FA fa_2310(.A(stage4_c34_c_fa0), .B(stage4_c34_c_fa1), .C(stage4_c34_c_fa2), .So(stage5_c35_s_fa0), .Co(stage5_c35_c_fa0));
    FA fa_2311(.A(stage4_c34_c_ha0), .B(stage4_c35_s_fa0), .C(stage4_c35_s_fa1), .So(stage5_c35_s_fa1), .Co(stage5_c35_c_fa1));
    HA ha_149(.A(stage4_c35_s_fa2), .B(stage4_c35_s_ha0), .So(stage5_c35_s_ha0), .Co(stage5_c35_c_ha0));
    FA fa_2312(.A(stage4_c35_c_fa0), .B(stage4_c35_c_fa1), .C(stage4_c35_c_fa2), .So(stage5_c36_s_fa0), .Co(stage5_c36_c_fa0));
    FA fa_2313(.A(stage4_c35_c_ha0), .B(stage4_c36_s_fa0), .C(stage4_c36_s_fa1), .So(stage5_c36_s_fa1), .Co(stage5_c36_c_fa1));
    HA ha_150(.A(stage4_c36_s_fa2), .B(stage4_c36_s_ha0), .So(stage5_c36_s_ha0), .Co(stage5_c36_c_ha0));
    FA fa_2314(.A(stage4_c36_c_fa0), .B(stage4_c36_c_fa1), .C(stage4_c36_c_fa2), .So(stage5_c37_s_fa0), .Co(stage5_c37_c_fa0));
    FA fa_2315(.A(stage4_c36_c_ha0), .B(stage4_c37_s_fa0), .C(stage4_c37_s_fa1), .So(stage5_c37_s_fa1), .Co(stage5_c37_c_fa1));
    HA ha_151(.A(stage4_c37_s_fa2), .B(stage4_c37_s_fa3), .So(stage5_c37_s_ha0), .Co(stage5_c37_c_ha0));
    FA fa_2316(.A(stage4_c37_c_fa0), .B(stage4_c37_c_fa1), .C(stage4_c37_c_fa2), .So(stage5_c38_s_fa0), .Co(stage5_c38_c_fa0));
    FA fa_2317(.A(stage4_c37_c_fa3), .B(stage4_c38_s_fa0), .C(stage4_c38_s_fa1), .So(stage5_c38_s_fa1), .Co(stage5_c38_c_fa1));
    HA ha_152(.A(stage4_c38_s_fa2), .B(stage4_c38_s_fa3), .So(stage5_c38_s_ha0), .Co(stage5_c38_c_ha0));
    FA fa_2318(.A(stage4_c38_c_fa0), .B(stage4_c38_c_fa1), .C(stage4_c38_c_fa2), .So(stage5_c39_s_fa0), .Co(stage5_c39_c_fa0));
    FA fa_2319(.A(stage4_c38_c_fa3), .B(stage4_c39_s_fa0), .C(stage4_c39_s_fa1), .So(stage5_c39_s_fa1), .Co(stage5_c39_c_fa1));
    HA ha_153(.A(stage4_c39_s_fa2), .B(stage4_c39_s_fa3), .So(stage5_c39_s_ha0), .Co(stage5_c39_c_ha0));
    FA fa_2320(.A(stage4_c39_c_fa0), .B(stage4_c39_c_fa1), .C(stage4_c39_c_fa2), .So(stage5_c40_s_fa0), .Co(stage5_c40_c_fa0));
    FA fa_2321(.A(stage4_c39_c_fa3), .B(stage4_c40_s_fa0), .C(stage4_c40_s_fa1), .So(stage5_c40_s_fa1), .Co(stage5_c40_c_fa1));
    HA ha_154(.A(stage4_c40_s_fa2), .B(stage4_c40_s_fa3), .So(stage5_c40_s_ha0), .Co(stage5_c40_c_ha0));
    FA fa_2322(.A(stage4_c40_c_fa0), .B(stage4_c40_c_fa1), .C(stage4_c40_c_fa2), .So(stage5_c41_s_fa0), .Co(stage5_c41_c_fa0));
    FA fa_2323(.A(stage4_c40_c_fa3), .B(stage4_c41_s_fa0), .C(stage4_c41_s_fa1), .So(stage5_c41_s_fa1), .Co(stage5_c41_c_fa1));
    FA fa_2324(.A(stage4_c41_s_fa2), .B(stage4_c41_s_fa3), .C(stage1_c41_s_ha0), .So(stage5_c41_s_fa2), .Co(stage5_c41_c_fa2));
    FA fa_2325(.A(stage4_c41_c_fa0), .B(stage4_c41_c_fa1), .C(stage4_c41_c_fa2), .So(stage5_c42_s_fa0), .Co(stage5_c42_c_fa0));
    FA fa_2326(.A(stage4_c41_c_fa3), .B(stage4_c42_s_fa0), .C(stage4_c42_s_fa1), .So(stage5_c42_s_fa1), .Co(stage5_c42_c_fa1));
    FA fa_2327(.A(stage4_c42_s_fa2), .B(stage4_c42_s_fa3), .C(stage1_c42_s_ha0), .So(stage5_c42_s_fa2), .Co(stage5_c42_c_fa2));
    FA fa_2328(.A(stage4_c42_c_fa0), .B(stage4_c42_c_fa1), .C(stage4_c42_c_fa2), .So(stage5_c43_s_fa0), .Co(stage5_c43_c_fa0));
    FA fa_2329(.A(stage4_c42_c_fa3), .B(stage4_c43_s_fa0), .C(stage4_c43_s_fa1), .So(stage5_c43_s_fa1), .Co(stage5_c43_c_fa1));
    FA fa_2330(.A(stage4_c43_s_fa2), .B(stage4_c43_s_fa3), .C(stage1_c43_s_ha0), .So(stage5_c43_s_fa2), .Co(stage5_c43_c_fa2));
    FA fa_2331(.A(stage4_c43_c_fa0), .B(stage4_c43_c_fa1), .C(stage4_c43_c_fa2), .So(stage5_c44_s_fa0), .Co(stage5_c44_c_fa0));
    FA fa_2332(.A(stage4_c43_c_fa3), .B(stage4_c44_s_fa0), .C(stage4_c44_s_fa1), .So(stage5_c44_s_fa1), .Co(stage5_c44_c_fa1));
    FA fa_2333(.A(stage4_c44_s_fa2), .B(stage4_c44_s_fa3), .C(stage1_c44_s_ha0), .So(stage5_c44_s_fa2), .Co(stage5_c44_c_fa2));
    FA fa_2334(.A(stage4_c44_c_fa0), .B(stage4_c44_c_fa1), .C(stage4_c44_c_fa2), .So(stage5_c45_s_fa0), .Co(stage5_c45_c_fa0));
    FA fa_2335(.A(stage4_c44_c_fa3), .B(stage4_c45_s_fa0), .C(stage4_c45_s_fa1), .So(stage5_c45_s_fa1), .Co(stage5_c45_c_fa1));
    FA fa_2336(.A(stage4_c45_s_fa2), .B(stage4_c45_s_fa3), .C(stage1_c45_s_ha0), .So(stage5_c45_s_fa2), .Co(stage5_c45_c_fa2));
    FA fa_2337(.A(stage4_c45_c_fa0), .B(stage4_c45_c_fa1), .C(stage4_c45_c_fa2), .So(stage5_c46_s_fa0), .Co(stage5_c46_c_fa0));
    FA fa_2338(.A(stage4_c45_c_fa3), .B(stage4_c46_s_fa0), .C(stage4_c46_s_fa1), .So(stage5_c46_s_fa1), .Co(stage5_c46_c_fa1));
    FA fa_2339(.A(stage4_c46_s_fa2), .B(stage4_c46_s_fa3), .C(stage1_c46_s_ha0), .So(stage5_c46_s_fa2), .Co(stage5_c46_c_fa2));
    FA fa_2340(.A(stage4_c46_c_fa0), .B(stage4_c46_c_fa1), .C(stage4_c46_c_fa2), .So(stage5_c47_s_fa0), .Co(stage5_c47_c_fa0));
    FA fa_2341(.A(stage4_c46_c_fa3), .B(stage4_c47_s_fa0), .C(stage4_c47_s_fa1), .So(stage5_c47_s_fa1), .Co(stage5_c47_c_fa1));
    FA fa_2342(.A(stage4_c47_s_fa2), .B(stage4_c47_s_fa3), .C(stage1_c47_s_ha0), .So(stage5_c47_s_fa2), .Co(stage5_c47_c_fa2));
    FA fa_2343(.A(stage4_c47_c_fa0), .B(stage4_c47_c_fa1), .C(stage4_c47_c_fa2), .So(stage5_c48_s_fa0), .Co(stage5_c48_c_fa0));
    FA fa_2344(.A(stage4_c47_c_fa3), .B(stage4_c48_s_fa0), .C(stage4_c48_s_fa1), .So(stage5_c48_s_fa1), .Co(stage5_c48_c_fa1));
    FA fa_2345(.A(stage4_c48_s_fa2), .B(stage4_c48_s_fa3), .C(stage1_c48_s_ha0), .So(stage5_c48_s_fa2), .Co(stage5_c48_c_fa2));
    FA fa_2346(.A(stage4_c48_c_fa0), .B(stage4_c48_c_fa1), .C(stage4_c48_c_fa2), .So(stage5_c49_s_fa0), .Co(stage5_c49_c_fa0));
    FA fa_2347(.A(stage4_c48_c_fa3), .B(stage4_c49_s_fa0), .C(stage4_c49_s_fa1), .So(stage5_c49_s_fa1), .Co(stage5_c49_c_fa1));
    FA fa_2348(.A(stage4_c49_s_fa2), .B(stage4_c49_s_fa3), .C(stage1_c49_s_ha0), .So(stage5_c49_s_fa2), .Co(stage5_c49_c_fa2));
    FA fa_2349(.A(stage4_c49_c_fa0), .B(stage4_c49_c_fa1), .C(stage4_c49_c_fa2), .So(stage5_c50_s_fa0), .Co(stage5_c50_c_fa0));
    FA fa_2350(.A(stage4_c49_c_fa3), .B(stage4_c50_s_fa0), .C(stage4_c50_s_fa1), .So(stage5_c50_s_fa1), .Co(stage5_c50_c_fa1));
    FA fa_2351(.A(stage4_c50_s_fa2), .B(stage4_c50_s_fa3), .C(stage1_c50_s_ha0), .So(stage5_c50_s_fa2), .Co(stage5_c50_c_fa2));
    FA fa_2352(.A(stage4_c50_c_fa0), .B(stage4_c50_c_fa1), .C(stage4_c50_c_fa2), .So(stage5_c51_s_fa0), .Co(stage5_c51_c_fa0));
    FA fa_2353(.A(stage4_c50_c_fa3), .B(stage4_c51_s_fa0), .C(stage4_c51_s_fa1), .So(stage5_c51_s_fa1), .Co(stage5_c51_c_fa1));
    FA fa_2354(.A(stage4_c51_s_fa2), .B(stage4_c51_s_fa3), .C(stage1_c51_s_ha0), .So(stage5_c51_s_fa2), .Co(stage5_c51_c_fa2));
    FA fa_2355(.A(stage4_c51_c_fa0), .B(stage4_c51_c_fa1), .C(stage4_c51_c_fa2), .So(stage5_c52_s_fa0), .Co(stage5_c52_c_fa0));
    FA fa_2356(.A(stage4_c51_c_fa3), .B(stage4_c52_s_fa0), .C(stage4_c52_s_fa1), .So(stage5_c52_s_fa1), .Co(stage5_c52_c_fa1));
    FA fa_2357(.A(stage4_c52_s_fa2), .B(stage4_c52_s_fa3), .C(stage1_c52_s_ha0), .So(stage5_c52_s_fa2), .Co(stage5_c52_c_fa2));
    FA fa_2358(.A(stage4_c52_c_fa0), .B(stage4_c52_c_fa1), .C(stage4_c52_c_fa2), .So(stage5_c53_s_fa0), .Co(stage5_c53_c_fa0));
    FA fa_2359(.A(stage4_c52_c_fa3), .B(stage4_c53_s_fa0), .C(stage4_c53_s_fa1), .So(stage5_c53_s_fa1), .Co(stage5_c53_c_fa1));
    FA fa_2360(.A(stage4_c53_s_fa2), .B(stage4_c53_s_fa3), .C(stage1_c53_s_ha0), .So(stage5_c53_s_fa2), .Co(stage5_c53_c_fa2));
    FA fa_2361(.A(stage4_c53_c_fa0), .B(stage4_c53_c_fa1), .C(stage4_c53_c_fa2), .So(stage5_c54_s_fa0), .Co(stage5_c54_c_fa0));
    FA fa_2362(.A(stage4_c53_c_fa3), .B(stage4_c54_s_fa0), .C(stage4_c54_s_fa1), .So(stage5_c54_s_fa1), .Co(stage5_c54_c_fa1));
    FA fa_2363(.A(stage4_c54_s_fa2), .B(stage4_c54_s_fa3), .C(stage1_c54_s_ha0), .So(stage5_c54_s_fa2), .Co(stage5_c54_c_fa2));
    FA fa_2364(.A(stage4_c54_c_fa0), .B(stage4_c54_c_fa1), .C(stage4_c54_c_fa2), .So(stage5_c55_s_fa0), .Co(stage5_c55_c_fa0));
    FA fa_2365(.A(stage4_c54_c_fa3), .B(stage4_c55_s_fa0), .C(stage4_c55_s_fa1), .So(stage5_c55_s_fa1), .Co(stage5_c55_c_fa1));
    FA fa_2366(.A(stage4_c55_s_fa2), .B(stage4_c55_s_fa3), .C(stage1_c55_s_ha0), .So(stage5_c55_s_fa2), .Co(stage5_c55_c_fa2));
    FA fa_2367(.A(stage4_c55_c_fa0), .B(stage4_c55_c_fa1), .C(stage4_c55_c_fa2), .So(stage5_c56_s_fa0), .Co(stage5_c56_c_fa0));
    FA fa_2368(.A(stage4_c55_c_fa3), .B(stage4_c56_s_fa0), .C(stage4_c56_s_fa1), .So(stage5_c56_s_fa1), .Co(stage5_c56_c_fa1));
    FA fa_2369(.A(stage4_c56_s_fa2), .B(stage4_c56_s_fa3), .C(stage1_c56_s_ha0), .So(stage5_c56_s_fa2), .Co(stage5_c56_c_fa2));
    FA fa_2370(.A(stage4_c56_c_fa0), .B(stage4_c56_c_fa1), .C(stage4_c56_c_fa2), .So(stage5_c57_s_fa0), .Co(stage5_c57_c_fa0));
    FA fa_2371(.A(stage4_c56_c_fa3), .B(stage4_c57_s_fa0), .C(stage4_c57_s_fa1), .So(stage5_c57_s_fa1), .Co(stage5_c57_c_fa1));
    FA fa_2372(.A(stage4_c57_s_fa2), .B(stage4_c57_s_fa3), .C(stage1_c57_s_ha0), .So(stage5_c57_s_fa2), .Co(stage5_c57_c_fa2));
    FA fa_2373(.A(stage4_c57_c_fa0), .B(stage4_c57_c_fa1), .C(stage4_c57_c_fa2), .So(stage5_c58_s_fa0), .Co(stage5_c58_c_fa0));
    FA fa_2374(.A(stage4_c57_c_fa3), .B(stage4_c58_s_fa0), .C(stage4_c58_s_fa1), .So(stage5_c58_s_fa1), .Co(stage5_c58_c_fa1));
    FA fa_2375(.A(stage4_c58_s_fa2), .B(stage4_c58_s_fa3), .C(stage1_c58_s_ha0), .So(stage5_c58_s_fa2), .Co(stage5_c58_c_fa2));
    FA fa_2376(.A(stage4_c58_c_fa0), .B(stage4_c58_c_fa1), .C(stage4_c58_c_fa2), .So(stage5_c59_s_fa0), .Co(stage5_c59_c_fa0));
    FA fa_2377(.A(stage4_c58_c_fa3), .B(stage4_c59_s_fa0), .C(stage4_c59_s_fa1), .So(stage5_c59_s_fa1), .Co(stage5_c59_c_fa1));
    FA fa_2378(.A(stage4_c59_s_fa2), .B(stage4_c59_s_fa3), .C(stage1_c59_s_ha0), .So(stage5_c59_s_fa2), .Co(stage5_c59_c_fa2));
    FA fa_2379(.A(stage4_c59_c_fa0), .B(stage4_c59_c_fa1), .C(stage4_c59_c_fa2), .So(stage5_c60_s_fa0), .Co(stage5_c60_c_fa0));
    FA fa_2380(.A(stage4_c59_c_fa3), .B(stage4_c60_s_fa0), .C(stage4_c60_s_fa1), .So(stage5_c60_s_fa1), .Co(stage5_c60_c_fa1));
    FA fa_2381(.A(stage4_c60_s_fa2), .B(stage4_c60_s_fa3), .C(stage1_c60_s_ha0), .So(stage5_c60_s_fa2), .Co(stage5_c60_c_fa2));
    FA fa_2382(.A(stage4_c60_c_fa0), .B(stage4_c60_c_fa1), .C(stage4_c60_c_fa2), .So(stage5_c61_s_fa0), .Co(stage5_c61_c_fa0));
    FA fa_2383(.A(stage4_c60_c_fa3), .B(stage4_c61_s_fa0), .C(stage4_c61_s_fa1), .So(stage5_c61_s_fa1), .Co(stage5_c61_c_fa1));
    FA fa_2384(.A(stage4_c61_s_fa2), .B(stage4_c61_s_fa3), .C(stage1_c61_s_ha0), .So(stage5_c61_s_fa2), .Co(stage5_c61_c_fa2));
    FA fa_2385(.A(stage4_c61_c_fa0), .B(stage4_c61_c_fa1), .C(stage4_c61_c_fa2), .So(stage5_c62_s_fa0), .Co(stage5_c62_c_fa0));
    FA fa_2386(.A(stage4_c61_c_fa3), .B(stage4_c62_s_fa0), .C(stage4_c62_s_fa1), .So(stage5_c62_s_fa1), .Co(stage5_c62_c_fa1));
    FA fa_2387(.A(stage4_c62_s_fa2), .B(stage4_c62_s_fa3), .C(stage1_c62_s_ha0), .So(stage5_c62_s_fa2), .Co(stage5_c62_c_fa2));
    FA fa_2388(.A(stage4_c62_c_fa0), .B(stage4_c62_c_fa1), .C(stage4_c62_c_fa2), .So(stage5_c63_s_fa0), .Co(stage5_c63_c_fa0));
    FA fa_2389(.A(stage4_c62_c_fa3), .B(stage4_c63_s_fa0), .C(stage4_c63_s_fa1), .So(stage5_c63_s_fa1), .Co(stage5_c63_c_fa1));
    FA fa_2390(.A(stage4_c63_s_fa2), .B(stage4_c63_s_fa3), .C(stage1_c63_s_ha0), .So(stage5_c63_s_fa2), .Co(stage5_c63_c_fa2));
    FA fa_2391(.A(stage4_c63_c_fa0), .B(stage4_c63_c_fa1), .C(stage4_c63_c_fa2), .So(stage5_c64_s_fa0), .Co(stage5_c64_c_fa0));
    FA fa_2392(.A(stage4_c63_c_fa3), .B(stage4_c64_s_fa0), .C(stage4_c64_s_fa1), .So(stage5_c64_s_fa1), .Co(stage5_c64_c_fa1));
    FA fa_2393(.A(stage4_c64_s_fa2), .B(stage4_c64_s_fa3), .C(stage1_c64_s_ha0), .So(stage5_c64_s_fa2), .Co(stage5_c64_c_fa2));
    FA fa_2394(.A(stage4_c64_c_fa0), .B(stage4_c64_c_fa1), .C(stage4_c64_c_fa2), .So(stage5_c65_s_fa0), .Co(stage5_c65_c_fa0));
    FA fa_2395(.A(stage4_c64_c_fa3), .B(stage4_c65_s_fa0), .C(stage4_c65_s_fa1), .So(stage5_c65_s_fa1), .Co(stage5_c65_c_fa1));
    FA fa_2396(.A(stage4_c65_s_fa2), .B(stage4_c65_s_fa3), .C(stage1_c65_s_ha0), .So(stage5_c65_s_fa2), .Co(stage5_c65_c_fa2));
    FA fa_2397(.A(stage4_c65_c_fa0), .B(stage4_c65_c_fa1), .C(stage4_c65_c_fa2), .So(stage5_c66_s_fa0), .Co(stage5_c66_c_fa0));
    FA fa_2398(.A(stage4_c65_c_fa3), .B(stage4_c66_s_fa0), .C(stage4_c66_s_fa1), .So(stage5_c66_s_fa1), .Co(stage5_c66_c_fa1));
    FA fa_2399(.A(stage4_c66_s_fa2), .B(stage4_c66_s_fa3), .C(stage1_c66_s_ha0), .So(stage5_c66_s_fa2), .Co(stage5_c66_c_fa2));
    FA fa_2400(.A(stage4_c66_c_fa0), .B(stage4_c66_c_fa1), .C(stage4_c66_c_fa2), .So(stage5_c67_s_fa0), .Co(stage5_c67_c_fa0));
    FA fa_2401(.A(stage4_c66_c_fa3), .B(stage4_c67_s_fa0), .C(stage4_c67_s_fa1), .So(stage5_c67_s_fa1), .Co(stage5_c67_c_fa1));
    FA fa_2402(.A(stage4_c67_s_fa2), .B(stage4_c67_s_fa3), .C(stage1_c67_s_ha0), .So(stage5_c67_s_fa2), .Co(stage5_c67_c_fa2));
    FA fa_2403(.A(stage4_c67_c_fa0), .B(stage4_c67_c_fa1), .C(stage4_c67_c_fa2), .So(stage5_c68_s_fa0), .Co(stage5_c68_c_fa0));
    FA fa_2404(.A(stage4_c67_c_fa3), .B(stage4_c68_s_fa0), .C(stage4_c68_s_fa1), .So(stage5_c68_s_fa1), .Co(stage5_c68_c_fa1));
    FA fa_2405(.A(stage4_c68_s_fa2), .B(stage4_c68_s_fa3), .C(stage1_c68_s_ha0), .So(stage5_c68_s_fa2), .Co(stage5_c68_c_fa2));
    FA fa_2406(.A(stage4_c68_c_fa0), .B(stage4_c68_c_fa1), .C(stage4_c68_c_fa2), .So(stage5_c69_s_fa0), .Co(stage5_c69_c_fa0));
    FA fa_2407(.A(stage4_c68_c_fa3), .B(stage4_c69_s_fa0), .C(stage4_c69_s_fa1), .So(stage5_c69_s_fa1), .Co(stage5_c69_c_fa1));
    FA fa_2408(.A(stage4_c69_s_fa2), .B(stage4_c69_s_fa3), .C(stage1_c69_s_ha0), .So(stage5_c69_s_fa2), .Co(stage5_c69_c_fa2));
    FA fa_2409(.A(stage4_c69_c_fa0), .B(stage4_c69_c_fa1), .C(stage4_c69_c_fa2), .So(stage5_c70_s_fa0), .Co(stage5_c70_c_fa0));
    FA fa_2410(.A(stage4_c69_c_fa3), .B(stage4_c70_s_fa0), .C(stage4_c70_s_fa1), .So(stage5_c70_s_fa1), .Co(stage5_c70_c_fa1));
    FA fa_2411(.A(stage4_c70_s_fa2), .B(stage4_c70_s_fa3), .C(stage1_c70_s_ha0), .So(stage5_c70_s_fa2), .Co(stage5_c70_c_fa2));
    FA fa_2412(.A(stage4_c70_c_fa0), .B(stage4_c70_c_fa1), .C(stage4_c70_c_fa2), .So(stage5_c71_s_fa0), .Co(stage5_c71_c_fa0));
    FA fa_2413(.A(stage4_c70_c_fa3), .B(stage4_c71_s_fa0), .C(stage4_c71_s_fa1), .So(stage5_c71_s_fa1), .Co(stage5_c71_c_fa1));
    FA fa_2414(.A(stage4_c71_s_fa2), .B(stage4_c71_s_fa3), .C(stage1_c71_s_ha0), .So(stage5_c71_s_fa2), .Co(stage5_c71_c_fa2));
    FA fa_2415(.A(stage4_c71_c_fa0), .B(stage4_c71_c_fa1), .C(stage4_c71_c_fa2), .So(stage5_c72_s_fa0), .Co(stage5_c72_c_fa0));
    FA fa_2416(.A(stage4_c71_c_fa3), .B(stage4_c72_s_fa0), .C(stage4_c72_s_fa1), .So(stage5_c72_s_fa1), .Co(stage5_c72_c_fa1));
    FA fa_2417(.A(stage4_c72_s_fa2), .B(stage4_c72_s_fa3), .C(stage0_r71_c1), .So(stage5_c72_s_fa2), .Co(stage5_c72_c_fa2));
    FA fa_2418(.A(stage4_c72_c_fa0), .B(stage4_c72_c_fa1), .C(stage4_c72_c_fa2), .So(stage5_c73_s_fa0), .Co(stage5_c73_c_fa0));
    FA fa_2419(.A(stage4_c72_c_fa3), .B(stage4_c73_s_fa0), .C(stage4_c73_s_fa1), .So(stage5_c73_s_fa1), .Co(stage5_c73_c_fa1));
    HA ha_155(.A(stage4_c73_s_fa2), .B(stage4_c73_s_fa3), .So(stage5_c73_s_ha0), .Co(stage5_c73_c_ha0));
    FA fa_2420(.A(stage4_c73_c_fa0), .B(stage4_c73_c_fa1), .C(stage4_c73_c_fa2), .So(stage5_c74_s_fa0), .Co(stage5_c74_c_fa0));
    FA fa_2421(.A(stage4_c73_c_fa3), .B(stage4_c74_s_fa0), .C(stage4_c74_s_fa1), .So(stage5_c74_s_fa1), .Co(stage5_c74_c_fa1));
    HA ha_156(.A(stage4_c74_s_fa2), .B(stage4_c74_s_fa3), .So(stage5_c74_s_ha0), .Co(stage5_c74_c_ha0));
    FA fa_2422(.A(stage4_c74_c_fa0), .B(stage4_c74_c_fa1), .C(stage4_c74_c_fa2), .So(stage5_c75_s_fa0), .Co(stage5_c75_c_fa0));
    FA fa_2423(.A(stage4_c74_c_fa3), .B(stage4_c75_s_fa0), .C(stage4_c75_s_fa1), .So(stage5_c75_s_fa1), .Co(stage5_c75_c_fa1));
    HA ha_157(.A(stage4_c75_s_fa2), .B(stage4_c75_s_fa3), .So(stage5_c75_s_ha0), .Co(stage5_c75_c_ha0));
    FA fa_2424(.A(stage4_c75_c_fa0), .B(stage4_c75_c_fa1), .C(stage4_c75_c_fa2), .So(stage5_c76_s_fa0), .Co(stage5_c76_c_fa0));
    FA fa_2425(.A(stage4_c75_c_fa3), .B(stage4_c76_s_fa0), .C(stage4_c76_s_fa1), .So(stage5_c76_s_fa1), .Co(stage5_c76_c_fa1));
    HA ha_158(.A(stage4_c76_s_fa2), .B(stage4_c76_s_fa3), .So(stage5_c76_s_ha0), .Co(stage5_c76_c_ha0));
    FA fa_2426(.A(stage4_c76_c_fa0), .B(stage4_c76_c_fa1), .C(stage4_c76_c_fa2), .So(stage5_c77_s_fa0), .Co(stage5_c77_c_fa0));
    FA fa_2427(.A(stage4_c76_c_fa3), .B(stage4_c77_s_fa0), .C(stage4_c77_s_fa1), .So(stage5_c77_s_fa1), .Co(stage5_c77_c_fa1));
    HA ha_159(.A(stage4_c77_s_fa2), .B(stage4_c77_s_fa3), .So(stage5_c77_s_ha0), .Co(stage5_c77_c_ha0));
    FA fa_2428(.A(stage4_c77_c_fa0), .B(stage4_c77_c_fa1), .C(stage4_c77_c_fa2), .So(stage5_c78_s_fa0), .Co(stage5_c78_c_fa0));
    FA fa_2429(.A(stage4_c77_c_fa3), .B(stage4_c78_s_fa0), .C(stage4_c78_s_fa1), .So(stage5_c78_s_fa1), .Co(stage5_c78_c_fa1));
    HA ha_160(.A(stage4_c78_s_fa2), .B(stage4_c78_s_ha0), .So(stage5_c78_s_ha0), .Co(stage5_c78_c_ha0));
    FA fa_2430(.A(stage4_c78_c_fa0), .B(stage4_c78_c_fa1), .C(stage4_c78_c_fa2), .So(stage5_c79_s_fa0), .Co(stage5_c79_c_fa0));
    FA fa_2431(.A(stage4_c78_c_ha0), .B(stage4_c79_s_fa0), .C(stage4_c79_s_fa1), .So(stage5_c79_s_fa1), .Co(stage5_c79_c_fa1));
    HA ha_161(.A(stage4_c79_s_fa2), .B(stage4_c79_s_ha0), .So(stage5_c79_s_ha0), .Co(stage5_c79_c_ha0));
    FA fa_2432(.A(stage4_c79_c_fa0), .B(stage4_c79_c_fa1), .C(stage4_c79_c_fa2), .So(stage5_c80_s_fa0), .Co(stage5_c80_c_fa0));
    FA fa_2433(.A(stage4_c79_c_ha0), .B(stage4_c80_s_fa0), .C(stage4_c80_s_fa1), .So(stage5_c80_s_fa1), .Co(stage5_c80_c_fa1));
    HA ha_162(.A(stage4_c80_s_fa2), .B(stage3_c80_s_fa4), .So(stage5_c80_s_ha0), .Co(stage5_c80_c_ha0));
    FA fa_2434(.A(stage4_c80_c_fa0), .B(stage4_c80_c_fa1), .C(stage4_c80_c_fa2), .So(stage5_c81_s_fa0), .Co(stage5_c81_c_fa0));
    FA fa_2435(.A(stage4_c81_s_fa0), .B(stage4_c81_s_fa1), .C(stage4_c81_s_fa2), .So(stage5_c81_s_fa1), .Co(stage5_c81_c_fa1));
    FA fa_2436(.A(stage4_c81_c_fa0), .B(stage4_c81_c_fa1), .C(stage4_c81_c_fa2), .So(stage5_c82_s_fa0), .Co(stage5_c82_c_fa0));
    FA fa_2437(.A(stage4_c82_s_fa0), .B(stage4_c82_s_fa1), .C(stage4_c82_s_fa2), .So(stage5_c82_s_fa1), .Co(stage5_c82_c_fa1));
    FA fa_2438(.A(stage4_c82_c_fa0), .B(stage4_c82_c_fa1), .C(stage4_c82_c_fa2), .So(stage5_c83_s_fa0), .Co(stage5_c83_c_fa0));
    FA fa_2439(.A(stage4_c83_s_fa0), .B(stage4_c83_s_fa1), .C(stage4_c83_s_fa2), .So(stage5_c83_s_fa1), .Co(stage5_c83_c_fa1));
    FA fa_2440(.A(stage4_c83_c_fa0), .B(stage4_c83_c_fa1), .C(stage4_c83_c_fa2), .So(stage5_c84_s_fa0), .Co(stage5_c84_c_fa0));
    FA fa_2441(.A(stage4_c84_s_fa0), .B(stage4_c84_s_fa1), .C(stage4_c84_s_fa2), .So(stage5_c84_s_fa1), .Co(stage5_c84_c_fa1));
    FA fa_2442(.A(stage4_c84_c_fa0), .B(stage4_c84_c_fa1), .C(stage4_c84_c_fa2), .So(stage5_c85_s_fa0), .Co(stage5_c85_c_fa0));
    FA fa_2443(.A(stage4_c85_s_fa0), .B(stage4_c85_s_fa1), .C(stage4_c85_s_fa2), .So(stage5_c85_s_fa1), .Co(stage5_c85_c_fa1));
    FA fa_2444(.A(stage4_c85_c_fa0), .B(stage4_c85_c_fa1), .C(stage4_c85_c_fa2), .So(stage5_c86_s_fa0), .Co(stage5_c86_c_fa0));
    FA fa_2445(.A(stage4_c86_s_fa0), .B(stage4_c86_s_fa1), .C(stage4_c86_s_ha0), .So(stage5_c86_s_fa1), .Co(stage5_c86_c_fa1));
    FA fa_2446(.A(stage4_c86_c_fa0), .B(stage4_c86_c_fa1), .C(stage4_c86_c_ha0), .So(stage5_c87_s_fa0), .Co(stage5_c87_c_fa0));
    FA fa_2447(.A(stage4_c87_s_fa0), .B(stage4_c87_s_fa1), .C(stage4_c87_s_ha0), .So(stage5_c87_s_fa1), .Co(stage5_c87_c_fa1));
    FA fa_2448(.A(stage4_c87_c_fa0), .B(stage4_c87_c_fa1), .C(stage4_c87_c_ha0), .So(stage5_c88_s_fa0), .Co(stage5_c88_c_fa0));
    FA fa_2449(.A(stage4_c88_s_fa0), .B(stage4_c88_s_fa1), .C(stage4_c88_s_ha0), .So(stage5_c88_s_fa1), .Co(stage5_c88_c_fa1));
    FA fa_2450(.A(stage4_c88_c_fa0), .B(stage4_c88_c_fa1), .C(stage4_c88_c_ha0), .So(stage5_c89_s_fa0), .Co(stage5_c89_c_fa0));
    FA fa_2451(.A(stage4_c89_s_fa0), .B(stage4_c89_s_fa1), .C(stage4_c89_s_ha0), .So(stage5_c89_s_fa1), .Co(stage5_c89_c_fa1));
    FA fa_2452(.A(stage4_c89_c_fa0), .B(stage4_c89_c_fa1), .C(stage4_c89_c_ha0), .So(stage5_c90_s_fa0), .Co(stage5_c90_c_fa0));
    FA fa_2453(.A(stage4_c90_s_fa0), .B(stage4_c90_s_fa1), .C(stage4_c90_s_ha0), .So(stage5_c90_s_fa1), .Co(stage5_c90_c_fa1));
    FA fa_2454(.A(stage4_c90_c_fa0), .B(stage4_c90_c_fa1), .C(stage4_c90_c_ha0), .So(stage5_c91_s_fa0), .Co(stage5_c91_c_fa0));
    FA fa_2455(.A(stage4_c91_s_fa0), .B(stage4_c91_s_fa1), .C(stage4_c91_s_ha0), .So(stage5_c91_s_fa1), .Co(stage5_c91_c_fa1));
    FA fa_2456(.A(stage4_c91_c_fa0), .B(stage4_c91_c_fa1), .C(stage4_c91_c_ha0), .So(stage5_c92_s_fa0), .Co(stage5_c92_c_fa0));
    FA fa_2457(.A(stage4_c92_s_fa0), .B(stage4_c92_s_fa1), .C(stage2_c92_s_ha0), .So(stage5_c92_s_fa1), .Co(stage5_c92_c_fa1));
    FA fa_2458(.A(stage4_c92_c_fa0), .B(stage4_c92_c_fa1), .C(stage4_c93_s_fa0), .So(stage5_c93_s_fa0), .Co(stage5_c93_c_fa0));
    HA ha_163(.A(stage4_c93_s_fa1), .B(stage2_c93_s_ha0), .So(stage5_c93_s_ha0), .Co(stage5_c93_c_ha0));
    FA fa_2459(.A(stage4_c93_c_fa0), .B(stage4_c93_c_fa1), .C(stage4_c94_s_fa0), .So(stage5_c94_s_fa0), .Co(stage5_c94_c_fa0));
    FA fa_2460(.A(stage4_c94_c_fa0), .B(stage4_c94_c_fa1), .C(stage4_c95_s_fa0), .So(stage5_c95_s_fa0), .Co(stage5_c95_c_fa0));
    FA fa_2461(.A(stage4_c95_c_fa0), .B(stage4_c95_c_fa1), .C(stage4_c96_s_fa0), .So(stage5_c96_s_fa0), .Co(stage5_c96_c_fa0));
    FA fa_2462(.A(stage4_c96_c_fa0), .B(stage4_c96_c_fa1), .C(stage4_c97_s_fa0), .So(stage5_c97_s_fa0), .Co(stage5_c97_c_fa0));
    FA fa_2463(.A(stage4_c97_c_fa0), .B(stage4_c97_c_fa1), .C(stage4_c98_s_fa0), .So(stage5_c98_s_fa0), .Co(stage5_c98_c_fa0));
    FA fa_2464(.A(stage4_c98_c_fa0), .B(stage4_c98_c_fa1), .C(stage4_c99_s_fa0), .So(stage5_c99_s_fa0), .Co(stage5_c99_c_fa0));
    FA fa_2465(.A(stage4_c99_c_fa0), .B(stage4_c99_c_ha0), .C(stage4_c100_s_fa0), .So(stage5_c100_s_fa0), .Co(stage5_c100_c_fa0));
    FA fa_2466(.A(stage4_c100_c_fa0), .B(stage4_c101_s_fa0), .C(stage3_c101_s_fa1), .So(stage5_c101_s_fa0), .Co(stage5_c101_c_fa0));
    FA fa_2467(.A(stage4_c101_c_fa0), .B(stage4_c102_s_fa0), .C(stage3_c102_s_fa1), .So(stage5_c102_s_fa0), .Co(stage5_c102_c_fa0));
    FA fa_2468(.A(stage4_c102_c_fa0), .B(stage4_c103_s_fa0), .C(stage3_c103_s_ha0), .So(stage5_c103_s_fa0), .Co(stage5_c103_c_fa0));
    FA fa_2469(.A(stage4_c103_c_fa0), .B(stage4_c104_s_fa0), .C(stage2_c104_s_fa1), .So(stage5_c104_s_fa0), .Co(stage5_c104_c_fa0));
    HA ha_164(.A(stage4_c104_c_fa0), .B(stage4_c105_s_fa0), .So(stage5_c105_s_ha0), .Co(stage5_c105_c_ha0));
    HA ha_165(.A(stage4_c105_c_fa0), .B(stage4_c106_s_fa0), .So(stage5_c106_s_ha0), .Co(stage5_c106_c_ha0));
    HA ha_166(.A(stage4_c106_c_fa0), .B(stage4_c107_s_ha0), .So(stage5_c107_s_ha0), .Co(stage5_c107_c_ha0));
    HA ha_167(.A(stage4_c107_c_ha0), .B(stage4_c108_s_ha0), .So(stage5_c108_s_ha0), .Co(stage5_c108_c_ha0));
    HA ha_168(.A(stage4_c108_c_ha0), .B(stage4_c109_s_ha0), .So(stage5_c109_s_ha0), .Co(stage5_c109_c_ha0));
    HA ha_169(.A(stage4_c109_c_ha0), .B(stage4_c110_s_ha0), .So(stage5_c110_s_ha0), .Co(stage5_c110_c_ha0));
    HA ha_170(.A(stage4_c110_c_ha0), .B(stage4_c111_s_ha0), .So(stage5_c111_s_ha0), .Co(stage5_c111_c_ha0));
    HA ha_171(.A(stage4_c111_c_ha0), .B(stage4_c112_s_ha0), .So(stage5_c112_s_ha0), .Co(stage5_c112_c_ha0));
    HA ha_172(.A(stage5_c5_c_ha0), .B(stage5_c6_s_ha0), .So(stage6_c6_s_ha0), .Co(stage6_c6_c_ha0));
    HA ha_173(.A(stage5_c6_c_ha0), .B(stage5_c7_s_ha0), .So(stage6_c7_s_ha0), .Co(stage6_c7_c_ha0));
    HA ha_174(.A(stage5_c7_c_ha0), .B(stage5_c8_s_ha0), .So(stage6_c8_s_ha0), .Co(stage6_c8_c_ha0));
    HA ha_175(.A(stage5_c8_c_ha0), .B(stage5_c9_s_ha0), .So(stage6_c9_s_ha0), .Co(stage6_c9_c_ha0));
    HA ha_176(.A(stage5_c9_c_ha0), .B(stage5_c10_s_fa0), .So(stage6_c10_s_ha0), .Co(stage6_c10_c_ha0));
    HA ha_177(.A(stage5_c10_c_fa0), .B(stage5_c11_s_fa0), .So(stage6_c11_s_ha0), .Co(stage6_c11_c_ha0));
    HA ha_178(.A(stage5_c11_c_fa0), .B(stage5_c12_s_fa0), .So(stage6_c12_s_ha0), .Co(stage6_c12_c_ha0));
    HA ha_179(.A(stage5_c12_c_fa0), .B(stage5_c13_s_fa0), .So(stage6_c13_s_ha0), .Co(stage6_c13_c_ha0));
    HA ha_180(.A(stage5_c13_c_fa0), .B(stage5_c14_s_fa0), .So(stage6_c14_s_ha0), .Co(stage6_c14_c_ha0));
    FA fa_2470(.A(stage5_c14_c_fa0), .B(stage5_c15_s_fa0), .C(stage4_c15_s_ha0), .So(stage6_c15_s_fa0), .Co(stage6_c15_c_fa0));
    FA fa_2471(.A(stage5_c15_c_fa0), .B(stage5_c16_s_fa0), .C(stage4_c16_s_ha0), .So(stage6_c16_s_fa0), .Co(stage6_c16_c_fa0));
    FA fa_2472(.A(stage5_c16_c_fa0), .B(stage5_c17_s_fa0), .C(stage4_c17_s_fa1), .So(stage6_c17_s_fa0), .Co(stage6_c17_c_fa0));
    FA fa_2473(.A(stage5_c17_c_fa0), .B(stage5_c18_s_fa0), .C(stage4_c18_s_fa1), .So(stage6_c18_s_fa0), .Co(stage6_c18_c_fa0));
    FA fa_2474(.A(stage5_c18_c_fa0), .B(stage5_c19_s_fa0), .C(stage4_c19_s_fa1), .So(stage6_c19_s_fa0), .Co(stage6_c19_c_fa0));
    FA fa_2475(.A(stage5_c19_c_fa0), .B(stage5_c20_s_fa0), .C(stage4_c20_s_fa1), .So(stage6_c20_s_fa0), .Co(stage6_c20_c_fa0));
    FA fa_2476(.A(stage5_c20_c_fa0), .B(stage5_c21_s_fa0), .C(stage5_c21_s_ha0), .So(stage6_c21_s_fa0), .Co(stage6_c21_c_fa0));
    FA fa_2477(.A(stage5_c21_c_fa0), .B(stage5_c21_c_ha0), .C(stage5_c22_s_fa0), .So(stage6_c22_s_fa0), .Co(stage6_c22_c_fa0));
    FA fa_2478(.A(stage5_c22_c_fa0), .B(stage5_c22_c_ha0), .C(stage5_c23_s_fa0), .So(stage6_c23_s_fa0), .Co(stage6_c23_c_fa0));
    FA fa_2479(.A(stage5_c23_c_fa0), .B(stage5_c23_c_ha0), .C(stage5_c24_s_fa0), .So(stage6_c24_s_fa0), .Co(stage6_c24_c_fa0));
    FA fa_2480(.A(stage5_c24_c_fa0), .B(stage5_c24_c_ha0), .C(stage5_c25_s_fa0), .So(stage6_c25_s_fa0), .Co(stage6_c25_c_fa0));
    FA fa_2481(.A(stage5_c25_c_fa0), .B(stage5_c25_c_fa1), .C(stage5_c26_s_fa0), .So(stage6_c26_s_fa0), .Co(stage6_c26_c_fa0));
    FA fa_2482(.A(stage5_c26_c_fa0), .B(stage5_c26_c_fa1), .C(stage5_c27_s_fa0), .So(stage6_c27_s_fa0), .Co(stage6_c27_c_fa0));
    FA fa_2483(.A(stage5_c27_c_fa0), .B(stage5_c27_c_fa1), .C(stage5_c28_s_fa0), .So(stage6_c28_s_fa0), .Co(stage6_c28_c_fa0));
    FA fa_2484(.A(stage5_c28_c_fa0), .B(stage5_c28_c_fa1), .C(stage5_c29_s_fa0), .So(stage6_c29_s_fa0), .Co(stage6_c29_c_fa0));
    FA fa_2485(.A(stage5_c29_c_fa0), .B(stage5_c29_c_fa1), .C(stage5_c30_s_fa0), .So(stage6_c30_s_fa0), .Co(stage6_c30_c_fa0));
    FA fa_2486(.A(stage5_c30_c_fa0), .B(stage5_c30_c_fa1), .C(stage5_c31_s_fa0), .So(stage6_c31_s_fa0), .Co(stage6_c31_c_fa0));
    HA ha_181(.A(stage5_c31_s_fa1), .B(stage3_c31_s_ha0), .So(stage6_c31_s_ha0), .Co(stage6_c31_c_ha0));
    FA fa_2487(.A(stage5_c31_c_fa0), .B(stage5_c31_c_fa1), .C(stage5_c32_s_fa0), .So(stage6_c32_s_fa0), .Co(stage6_c32_c_fa0));
    HA ha_182(.A(stage5_c32_s_fa1), .B(stage3_c32_s_fa4), .So(stage6_c32_s_ha0), .Co(stage6_c32_c_ha0));
    FA fa_2488(.A(stage5_c32_c_fa0), .B(stage5_c32_c_fa1), .C(stage5_c33_s_fa0), .So(stage6_c33_s_fa0), .Co(stage6_c33_c_fa0));
    HA ha_183(.A(stage5_c33_s_fa1), .B(stage3_c33_s_fa4), .So(stage6_c33_s_ha0), .Co(stage6_c33_c_ha0));
    FA fa_2489(.A(stage5_c33_c_fa0), .B(stage5_c33_c_fa1), .C(stage5_c34_s_fa0), .So(stage6_c34_s_fa0), .Co(stage6_c34_c_fa0));
    HA ha_184(.A(stage5_c34_s_fa1), .B(stage4_c34_s_ha0), .So(stage6_c34_s_ha0), .Co(stage6_c34_c_ha0));
    FA fa_2490(.A(stage5_c34_c_fa0), .B(stage5_c34_c_fa1), .C(stage5_c35_s_fa0), .So(stage6_c35_s_fa0), .Co(stage6_c35_c_fa0));
    HA ha_185(.A(stage5_c35_s_fa1), .B(stage5_c35_s_ha0), .So(stage6_c35_s_ha0), .Co(stage6_c35_c_ha0));
    FA fa_2491(.A(stage5_c35_c_fa0), .B(stage5_c35_c_fa1), .C(stage5_c35_c_ha0), .So(stage6_c36_s_fa0), .Co(stage6_c36_c_fa0));
    FA fa_2492(.A(stage5_c36_s_fa0), .B(stage5_c36_s_fa1), .C(stage5_c36_s_ha0), .So(stage6_c36_s_fa1), .Co(stage6_c36_c_fa1));
    FA fa_2493(.A(stage5_c36_c_fa0), .B(stage5_c36_c_fa1), .C(stage5_c36_c_ha0), .So(stage6_c37_s_fa0), .Co(stage6_c37_c_fa0));
    FA fa_2494(.A(stage5_c37_s_fa0), .B(stage5_c37_s_fa1), .C(stage5_c37_s_ha0), .So(stage6_c37_s_fa1), .Co(stage6_c37_c_fa1));
    FA fa_2495(.A(stage5_c37_c_fa0), .B(stage5_c37_c_fa1), .C(stage5_c37_c_ha0), .So(stage6_c38_s_fa0), .Co(stage6_c38_c_fa0));
    FA fa_2496(.A(stage5_c38_s_fa0), .B(stage5_c38_s_fa1), .C(stage5_c38_s_ha0), .So(stage6_c38_s_fa1), .Co(stage6_c38_c_fa1));
    FA fa_2497(.A(stage5_c38_c_fa0), .B(stage5_c38_c_fa1), .C(stage5_c38_c_ha0), .So(stage6_c39_s_fa0), .Co(stage6_c39_c_fa0));
    FA fa_2498(.A(stage5_c39_s_fa0), .B(stage5_c39_s_fa1), .C(stage5_c39_s_ha0), .So(stage6_c39_s_fa1), .Co(stage6_c39_c_fa1));
    FA fa_2499(.A(stage5_c39_c_fa0), .B(stage5_c39_c_fa1), .C(stage5_c39_c_ha0), .So(stage6_c40_s_fa0), .Co(stage6_c40_c_fa0));
    FA fa_2500(.A(stage5_c40_s_fa0), .B(stage5_c40_s_fa1), .C(stage5_c40_s_ha0), .So(stage6_c40_s_fa1), .Co(stage6_c40_c_fa1));
    FA fa_2501(.A(stage5_c40_c_fa0), .B(stage5_c40_c_fa1), .C(stage5_c40_c_ha0), .So(stage6_c41_s_fa0), .Co(stage6_c41_c_fa0));
    FA fa_2502(.A(stage5_c41_s_fa0), .B(stage5_c41_s_fa1), .C(stage5_c41_s_fa2), .So(stage6_c41_s_fa1), .Co(stage6_c41_c_fa1));
    FA fa_2503(.A(stage5_c41_c_fa0), .B(stage5_c41_c_fa1), .C(stage5_c41_c_fa2), .So(stage6_c42_s_fa0), .Co(stage6_c42_c_fa0));
    FA fa_2504(.A(stage5_c42_s_fa0), .B(stage5_c42_s_fa1), .C(stage5_c42_s_fa2), .So(stage6_c42_s_fa1), .Co(stage6_c42_c_fa1));
    FA fa_2505(.A(stage5_c42_c_fa0), .B(stage5_c42_c_fa1), .C(stage5_c42_c_fa2), .So(stage6_c43_s_fa0), .Co(stage6_c43_c_fa0));
    FA fa_2506(.A(stage5_c43_s_fa0), .B(stage5_c43_s_fa1), .C(stage5_c43_s_fa2), .So(stage6_c43_s_fa1), .Co(stage6_c43_c_fa1));
    FA fa_2507(.A(stage5_c43_c_fa0), .B(stage5_c43_c_fa1), .C(stage5_c43_c_fa2), .So(stage6_c44_s_fa0), .Co(stage6_c44_c_fa0));
    FA fa_2508(.A(stage5_c44_s_fa0), .B(stage5_c44_s_fa1), .C(stage5_c44_s_fa2), .So(stage6_c44_s_fa1), .Co(stage6_c44_c_fa1));
    FA fa_2509(.A(stage5_c44_c_fa0), .B(stage5_c44_c_fa1), .C(stage5_c44_c_fa2), .So(stage6_c45_s_fa0), .Co(stage6_c45_c_fa0));
    FA fa_2510(.A(stage5_c45_s_fa0), .B(stage5_c45_s_fa1), .C(stage5_c45_s_fa2), .So(stage6_c45_s_fa1), .Co(stage6_c45_c_fa1));
    FA fa_2511(.A(stage5_c45_c_fa0), .B(stage5_c45_c_fa1), .C(stage5_c45_c_fa2), .So(stage6_c46_s_fa0), .Co(stage6_c46_c_fa0));
    FA fa_2512(.A(stage5_c46_s_fa0), .B(stage5_c46_s_fa1), .C(stage5_c46_s_fa2), .So(stage6_c46_s_fa1), .Co(stage6_c46_c_fa1));
    FA fa_2513(.A(stage5_c46_c_fa0), .B(stage5_c46_c_fa1), .C(stage5_c46_c_fa2), .So(stage6_c47_s_fa0), .Co(stage6_c47_c_fa0));
    FA fa_2514(.A(stage5_c47_s_fa0), .B(stage5_c47_s_fa1), .C(stage5_c47_s_fa2), .So(stage6_c47_s_fa1), .Co(stage6_c47_c_fa1));
    FA fa_2515(.A(stage5_c47_c_fa0), .B(stage5_c47_c_fa1), .C(stage5_c47_c_fa2), .So(stage6_c48_s_fa0), .Co(stage6_c48_c_fa0));
    FA fa_2516(.A(stage5_c48_s_fa0), .B(stage5_c48_s_fa1), .C(stage5_c48_s_fa2), .So(stage6_c48_s_fa1), .Co(stage6_c48_c_fa1));
    FA fa_2517(.A(stage5_c48_c_fa0), .B(stage5_c48_c_fa1), .C(stage5_c48_c_fa2), .So(stage6_c49_s_fa0), .Co(stage6_c49_c_fa0));
    FA fa_2518(.A(stage5_c49_s_fa0), .B(stage5_c49_s_fa1), .C(stage5_c49_s_fa2), .So(stage6_c49_s_fa1), .Co(stage6_c49_c_fa1));
    FA fa_2519(.A(stage5_c49_c_fa0), .B(stage5_c49_c_fa1), .C(stage5_c49_c_fa2), .So(stage6_c50_s_fa0), .Co(stage6_c50_c_fa0));
    FA fa_2520(.A(stage5_c50_s_fa0), .B(stage5_c50_s_fa1), .C(stage5_c50_s_fa2), .So(stage6_c50_s_fa1), .Co(stage6_c50_c_fa1));
    FA fa_2521(.A(stage5_c50_c_fa0), .B(stage5_c50_c_fa1), .C(stage5_c50_c_fa2), .So(stage6_c51_s_fa0), .Co(stage6_c51_c_fa0));
    FA fa_2522(.A(stage5_c51_s_fa0), .B(stage5_c51_s_fa1), .C(stage5_c51_s_fa2), .So(stage6_c51_s_fa1), .Co(stage6_c51_c_fa1));
    FA fa_2523(.A(stage5_c51_c_fa0), .B(stage5_c51_c_fa1), .C(stage5_c51_c_fa2), .So(stage6_c52_s_fa0), .Co(stage6_c52_c_fa0));
    FA fa_2524(.A(stage5_c52_s_fa0), .B(stage5_c52_s_fa1), .C(stage5_c52_s_fa2), .So(stage6_c52_s_fa1), .Co(stage6_c52_c_fa1));
    FA fa_2525(.A(stage5_c52_c_fa0), .B(stage5_c52_c_fa1), .C(stage5_c52_c_fa2), .So(stage6_c53_s_fa0), .Co(stage6_c53_c_fa0));
    FA fa_2526(.A(stage5_c53_s_fa0), .B(stage5_c53_s_fa1), .C(stage5_c53_s_fa2), .So(stage6_c53_s_fa1), .Co(stage6_c53_c_fa1));
    FA fa_2527(.A(stage5_c53_c_fa0), .B(stage5_c53_c_fa1), .C(stage5_c53_c_fa2), .So(stage6_c54_s_fa0), .Co(stage6_c54_c_fa0));
    FA fa_2528(.A(stage5_c54_s_fa0), .B(stage5_c54_s_fa1), .C(stage5_c54_s_fa2), .So(stage6_c54_s_fa1), .Co(stage6_c54_c_fa1));
    FA fa_2529(.A(stage5_c54_c_fa0), .B(stage5_c54_c_fa1), .C(stage5_c54_c_fa2), .So(stage6_c55_s_fa0), .Co(stage6_c55_c_fa0));
    FA fa_2530(.A(stage5_c55_s_fa0), .B(stage5_c55_s_fa1), .C(stage5_c55_s_fa2), .So(stage6_c55_s_fa1), .Co(stage6_c55_c_fa1));
    FA fa_2531(.A(stage5_c55_c_fa0), .B(stage5_c55_c_fa1), .C(stage5_c55_c_fa2), .So(stage6_c56_s_fa0), .Co(stage6_c56_c_fa0));
    FA fa_2532(.A(stage5_c56_s_fa0), .B(stage5_c56_s_fa1), .C(stage5_c56_s_fa2), .So(stage6_c56_s_fa1), .Co(stage6_c56_c_fa1));
    FA fa_2533(.A(stage5_c56_c_fa0), .B(stage5_c56_c_fa1), .C(stage5_c56_c_fa2), .So(stage6_c57_s_fa0), .Co(stage6_c57_c_fa0));
    FA fa_2534(.A(stage5_c57_s_fa0), .B(stage5_c57_s_fa1), .C(stage5_c57_s_fa2), .So(stage6_c57_s_fa1), .Co(stage6_c57_c_fa1));
    FA fa_2535(.A(stage5_c57_c_fa0), .B(stage5_c57_c_fa1), .C(stage5_c57_c_fa2), .So(stage6_c58_s_fa0), .Co(stage6_c58_c_fa0));
    FA fa_2536(.A(stage5_c58_s_fa0), .B(stage5_c58_s_fa1), .C(stage5_c58_s_fa2), .So(stage6_c58_s_fa1), .Co(stage6_c58_c_fa1));
    FA fa_2537(.A(stage5_c58_c_fa0), .B(stage5_c58_c_fa1), .C(stage5_c58_c_fa2), .So(stage6_c59_s_fa0), .Co(stage6_c59_c_fa0));
    FA fa_2538(.A(stage5_c59_s_fa0), .B(stage5_c59_s_fa1), .C(stage5_c59_s_fa2), .So(stage6_c59_s_fa1), .Co(stage6_c59_c_fa1));
    FA fa_2539(.A(stage5_c59_c_fa0), .B(stage5_c59_c_fa1), .C(stage5_c59_c_fa2), .So(stage6_c60_s_fa0), .Co(stage6_c60_c_fa0));
    FA fa_2540(.A(stage5_c60_s_fa0), .B(stage5_c60_s_fa1), .C(stage5_c60_s_fa2), .So(stage6_c60_s_fa1), .Co(stage6_c60_c_fa1));
    FA fa_2541(.A(stage5_c60_c_fa0), .B(stage5_c60_c_fa1), .C(stage5_c60_c_fa2), .So(stage6_c61_s_fa0), .Co(stage6_c61_c_fa0));
    FA fa_2542(.A(stage5_c61_s_fa0), .B(stage5_c61_s_fa1), .C(stage5_c61_s_fa2), .So(stage6_c61_s_fa1), .Co(stage6_c61_c_fa1));
    FA fa_2543(.A(stage5_c61_c_fa0), .B(stage5_c61_c_fa1), .C(stage5_c61_c_fa2), .So(stage6_c62_s_fa0), .Co(stage6_c62_c_fa0));
    FA fa_2544(.A(stage5_c62_s_fa0), .B(stage5_c62_s_fa1), .C(stage5_c62_s_fa2), .So(stage6_c62_s_fa1), .Co(stage6_c62_c_fa1));
    FA fa_2545(.A(stage5_c62_c_fa0), .B(stage5_c62_c_fa1), .C(stage5_c62_c_fa2), .So(stage6_c63_s_fa0), .Co(stage6_c63_c_fa0));
    FA fa_2546(.A(stage5_c63_s_fa0), .B(stage5_c63_s_fa1), .C(stage5_c63_s_fa2), .So(stage6_c63_s_fa1), .Co(stage6_c63_c_fa1));
    FA fa_2547(.A(stage5_c63_c_fa0), .B(stage5_c63_c_fa1), .C(stage5_c63_c_fa2), .So(stage6_c64_s_fa0), .Co(stage6_c64_c_fa0));
    FA fa_2548(.A(stage5_c64_s_fa0), .B(stage5_c64_s_fa1), .C(stage5_c64_s_fa2), .So(stage6_c64_s_fa1), .Co(stage6_c64_c_fa1));
    FA fa_2549(.A(stage5_c64_c_fa0), .B(stage5_c64_c_fa1), .C(stage5_c64_c_fa2), .So(stage6_c65_s_fa0), .Co(stage6_c65_c_fa0));
    FA fa_2550(.A(stage5_c65_s_fa0), .B(stage5_c65_s_fa1), .C(stage5_c65_s_fa2), .So(stage6_c65_s_fa1), .Co(stage6_c65_c_fa1));
    FA fa_2551(.A(stage5_c65_c_fa0), .B(stage5_c65_c_fa1), .C(stage5_c65_c_fa2), .So(stage6_c66_s_fa0), .Co(stage6_c66_c_fa0));
    FA fa_2552(.A(stage5_c66_s_fa0), .B(stage5_c66_s_fa1), .C(stage5_c66_s_fa2), .So(stage6_c66_s_fa1), .Co(stage6_c66_c_fa1));
    FA fa_2553(.A(stage5_c66_c_fa0), .B(stage5_c66_c_fa1), .C(stage5_c66_c_fa2), .So(stage6_c67_s_fa0), .Co(stage6_c67_c_fa0));
    FA fa_2554(.A(stage5_c67_s_fa0), .B(stage5_c67_s_fa1), .C(stage5_c67_s_fa2), .So(stage6_c67_s_fa1), .Co(stage6_c67_c_fa1));
    FA fa_2555(.A(stage5_c67_c_fa0), .B(stage5_c67_c_fa1), .C(stage5_c67_c_fa2), .So(stage6_c68_s_fa0), .Co(stage6_c68_c_fa0));
    FA fa_2556(.A(stage5_c68_s_fa0), .B(stage5_c68_s_fa1), .C(stage5_c68_s_fa2), .So(stage6_c68_s_fa1), .Co(stage6_c68_c_fa1));
    FA fa_2557(.A(stage5_c68_c_fa0), .B(stage5_c68_c_fa1), .C(stage5_c68_c_fa2), .So(stage6_c69_s_fa0), .Co(stage6_c69_c_fa0));
    FA fa_2558(.A(stage5_c69_s_fa0), .B(stage5_c69_s_fa1), .C(stage5_c69_s_fa2), .So(stage6_c69_s_fa1), .Co(stage6_c69_c_fa1));
    FA fa_2559(.A(stage5_c69_c_fa0), .B(stage5_c69_c_fa1), .C(stage5_c69_c_fa2), .So(stage6_c70_s_fa0), .Co(stage6_c70_c_fa0));
    FA fa_2560(.A(stage5_c70_s_fa0), .B(stage5_c70_s_fa1), .C(stage5_c70_s_fa2), .So(stage6_c70_s_fa1), .Co(stage6_c70_c_fa1));
    FA fa_2561(.A(stage5_c70_c_fa0), .B(stage5_c70_c_fa1), .C(stage5_c70_c_fa2), .So(stage6_c71_s_fa0), .Co(stage6_c71_c_fa0));
    FA fa_2562(.A(stage5_c71_s_fa0), .B(stage5_c71_s_fa1), .C(stage5_c71_s_fa2), .So(stage6_c71_s_fa1), .Co(stage6_c71_c_fa1));
    FA fa_2563(.A(stage5_c71_c_fa0), .B(stage5_c71_c_fa1), .C(stage5_c71_c_fa2), .So(stage6_c72_s_fa0), .Co(stage6_c72_c_fa0));
    FA fa_2564(.A(stage5_c72_s_fa0), .B(stage5_c72_s_fa1), .C(stage5_c72_s_fa2), .So(stage6_c72_s_fa1), .Co(stage6_c72_c_fa1));
    FA fa_2565(.A(stage5_c72_c_fa0), .B(stage5_c72_c_fa1), .C(stage5_c72_c_fa2), .So(stage6_c73_s_fa0), .Co(stage6_c73_c_fa0));
    FA fa_2566(.A(stage5_c73_s_fa0), .B(stage5_c73_s_fa1), .C(stage5_c73_s_ha0), .So(stage6_c73_s_fa1), .Co(stage6_c73_c_fa1));
    FA fa_2567(.A(stage5_c73_c_fa0), .B(stage5_c73_c_fa1), .C(stage5_c73_c_ha0), .So(stage6_c74_s_fa0), .Co(stage6_c74_c_fa0));
    FA fa_2568(.A(stage5_c74_s_fa0), .B(stage5_c74_s_fa1), .C(stage5_c74_s_ha0), .So(stage6_c74_s_fa1), .Co(stage6_c74_c_fa1));
    FA fa_2569(.A(stage5_c74_c_fa0), .B(stage5_c74_c_fa1), .C(stage5_c74_c_ha0), .So(stage6_c75_s_fa0), .Co(stage6_c75_c_fa0));
    FA fa_2570(.A(stage5_c75_s_fa0), .B(stage5_c75_s_fa1), .C(stage5_c75_s_ha0), .So(stage6_c75_s_fa1), .Co(stage6_c75_c_fa1));
    FA fa_2571(.A(stage5_c75_c_fa0), .B(stage5_c75_c_fa1), .C(stage5_c75_c_ha0), .So(stage6_c76_s_fa0), .Co(stage6_c76_c_fa0));
    FA fa_2572(.A(stage5_c76_s_fa0), .B(stage5_c76_s_fa1), .C(stage5_c76_s_ha0), .So(stage6_c76_s_fa1), .Co(stage6_c76_c_fa1));
    FA fa_2573(.A(stage5_c76_c_fa0), .B(stage5_c76_c_fa1), .C(stage5_c76_c_ha0), .So(stage6_c77_s_fa0), .Co(stage6_c77_c_fa0));
    FA fa_2574(.A(stage5_c77_s_fa0), .B(stage5_c77_s_fa1), .C(stage5_c77_s_ha0), .So(stage6_c77_s_fa1), .Co(stage6_c77_c_fa1));
    FA fa_2575(.A(stage5_c77_c_fa0), .B(stage5_c77_c_fa1), .C(stage5_c77_c_ha0), .So(stage6_c78_s_fa0), .Co(stage6_c78_c_fa0));
    FA fa_2576(.A(stage5_c78_s_fa0), .B(stage5_c78_s_fa1), .C(stage5_c78_s_ha0), .So(stage6_c78_s_fa1), .Co(stage6_c78_c_fa1));
    FA fa_2577(.A(stage5_c78_c_fa0), .B(stage5_c78_c_fa1), .C(stage5_c78_c_ha0), .So(stage6_c79_s_fa0), .Co(stage6_c79_c_fa0));
    FA fa_2578(.A(stage5_c79_s_fa0), .B(stage5_c79_s_fa1), .C(stage5_c79_s_ha0), .So(stage6_c79_s_fa1), .Co(stage6_c79_c_fa1));
    FA fa_2579(.A(stage5_c79_c_fa0), .B(stage5_c79_c_fa1), .C(stage5_c79_c_ha0), .So(stage6_c80_s_fa0), .Co(stage6_c80_c_fa0));
    FA fa_2580(.A(stage5_c80_s_fa0), .B(stage5_c80_s_fa1), .C(stage5_c80_s_ha0), .So(stage6_c80_s_fa1), .Co(stage6_c80_c_fa1));
    FA fa_2581(.A(stage5_c80_c_fa0), .B(stage5_c80_c_fa1), .C(stage5_c80_c_ha0), .So(stage6_c81_s_fa0), .Co(stage6_c81_c_fa0));
    FA fa_2582(.A(stage5_c81_s_fa0), .B(stage5_c81_s_fa1), .C(stage3_c81_s_fa4), .So(stage6_c81_s_fa1), .Co(stage6_c81_c_fa1));
    FA fa_2583(.A(stage5_c81_c_fa0), .B(stage5_c81_c_fa1), .C(stage5_c82_s_fa0), .So(stage6_c82_s_fa0), .Co(stage6_c82_c_fa0));
    HA ha_186(.A(stage5_c82_s_fa1), .B(stage3_c82_s_ha0), .So(stage6_c82_s_ha0), .Co(stage6_c82_c_ha0));
    FA fa_2584(.A(stage5_c82_c_fa0), .B(stage5_c82_c_fa1), .C(stage5_c83_s_fa0), .So(stage6_c83_s_fa0), .Co(stage6_c83_c_fa0));
    HA ha_187(.A(stage5_c83_s_fa1), .B(stage3_c83_s_ha0), .So(stage6_c83_s_ha0), .Co(stage6_c83_c_ha0));
    FA fa_2585(.A(stage5_c83_c_fa0), .B(stage5_c83_c_fa1), .C(stage5_c84_s_fa0), .So(stage6_c84_s_fa0), .Co(stage6_c84_c_fa0));
    HA ha_188(.A(stage5_c84_s_fa1), .B(stage3_c84_s_ha0), .So(stage6_c84_s_ha0), .Co(stage6_c84_c_ha0));
    FA fa_2586(.A(stage5_c84_c_fa0), .B(stage5_c84_c_fa1), .C(stage5_c85_s_fa0), .So(stage6_c85_s_fa0), .Co(stage6_c85_c_fa0));
    HA ha_189(.A(stage5_c85_s_fa1), .B(stage2_c85_s_fa5), .So(stage6_c85_s_ha0), .Co(stage6_c85_c_ha0));
    FA fa_2587(.A(stage5_c85_c_fa0), .B(stage5_c85_c_fa1), .C(stage5_c86_s_fa0), .So(stage6_c86_s_fa0), .Co(stage6_c86_c_fa0));
    FA fa_2588(.A(stage5_c86_c_fa0), .B(stage5_c86_c_fa1), .C(stage5_c87_s_fa0), .So(stage6_c87_s_fa0), .Co(stage6_c87_c_fa0));
    FA fa_2589(.A(stage5_c87_c_fa0), .B(stage5_c87_c_fa1), .C(stage5_c88_s_fa0), .So(stage6_c88_s_fa0), .Co(stage6_c88_c_fa0));
    FA fa_2590(.A(stage5_c88_c_fa0), .B(stage5_c88_c_fa1), .C(stage5_c89_s_fa0), .So(stage6_c89_s_fa0), .Co(stage6_c89_c_fa0));
    FA fa_2591(.A(stage5_c89_c_fa0), .B(stage5_c89_c_fa1), .C(stage5_c90_s_fa0), .So(stage6_c90_s_fa0), .Co(stage6_c90_c_fa0));
    FA fa_2592(.A(stage5_c90_c_fa0), .B(stage5_c90_c_fa1), .C(stage5_c91_s_fa0), .So(stage6_c91_s_fa0), .Co(stage6_c91_c_fa0));
    FA fa_2593(.A(stage5_c91_c_fa0), .B(stage5_c91_c_fa1), .C(stage5_c92_s_fa0), .So(stage6_c92_s_fa0), .Co(stage6_c92_c_fa0));
    FA fa_2594(.A(stage5_c92_c_fa0), .B(stage5_c92_c_fa1), .C(stage5_c93_s_fa0), .So(stage6_c93_s_fa0), .Co(stage6_c93_c_fa0));
    FA fa_2595(.A(stage5_c93_c_fa0), .B(stage5_c93_c_ha0), .C(stage5_c94_s_fa0), .So(stage6_c94_s_fa0), .Co(stage6_c94_c_fa0));
    FA fa_2596(.A(stage5_c94_c_fa0), .B(stage5_c95_s_fa0), .C(stage4_c95_s_fa1), .So(stage6_c95_s_fa0), .Co(stage6_c95_c_fa0));
    FA fa_2597(.A(stage5_c95_c_fa0), .B(stage5_c96_s_fa0), .C(stage4_c96_s_fa1), .So(stage6_c96_s_fa0), .Co(stage6_c96_c_fa0));
    FA fa_2598(.A(stage5_c96_c_fa0), .B(stage5_c97_s_fa0), .C(stage4_c97_s_fa1), .So(stage6_c97_s_fa0), .Co(stage6_c97_c_fa0));
    FA fa_2599(.A(stage5_c97_c_fa0), .B(stage5_c98_s_fa0), .C(stage4_c98_s_fa1), .So(stage6_c98_s_fa0), .Co(stage6_c98_c_fa0));
    FA fa_2600(.A(stage5_c98_c_fa0), .B(stage5_c99_s_fa0), .C(stage4_c99_s_ha0), .So(stage6_c99_s_fa0), .Co(stage6_c99_c_fa0));
    FA fa_2601(.A(stage5_c99_c_fa0), .B(stage5_c100_s_fa0), .C(stage3_c100_s_fa1), .So(stage6_c100_s_fa0), .Co(stage6_c100_c_fa0));
    HA ha_190(.A(stage5_c100_c_fa0), .B(stage5_c101_s_fa0), .So(stage6_c101_s_ha0), .Co(stage6_c101_c_ha0));
    HA ha_191(.A(stage5_c101_c_fa0), .B(stage5_c102_s_fa0), .So(stage6_c102_s_ha0), .Co(stage6_c102_c_ha0));
    HA ha_192(.A(stage5_c102_c_fa0), .B(stage5_c103_s_fa0), .So(stage6_c103_s_ha0), .Co(stage6_c103_c_ha0));
    HA ha_193(.A(stage5_c103_c_fa0), .B(stage5_c104_s_fa0), .So(stage6_c104_s_ha0), .Co(stage6_c104_c_ha0));
    HA ha_194(.A(stage5_c104_c_fa0), .B(stage5_c105_s_ha0), .So(stage6_c105_s_ha0), .Co(stage6_c105_c_ha0));
    HA ha_195(.A(stage5_c105_c_ha0), .B(stage5_c106_s_ha0), .So(stage6_c106_s_ha0), .Co(stage6_c106_c_ha0));
    HA ha_196(.A(stage5_c106_c_ha0), .B(stage5_c107_s_ha0), .So(stage6_c107_s_ha0), .Co(stage6_c107_c_ha0));
    HA ha_197(.A(stage5_c107_c_ha0), .B(stage5_c108_s_ha0), .So(stage6_c108_s_ha0), .Co(stage6_c108_c_ha0));
    HA ha_198(.A(stage5_c108_c_ha0), .B(stage5_c109_s_ha0), .So(stage6_c109_s_ha0), .Co(stage6_c109_c_ha0));
    HA ha_199(.A(stage5_c109_c_ha0), .B(stage5_c110_s_ha0), .So(stage6_c110_s_ha0), .Co(stage6_c110_c_ha0));
    HA ha_200(.A(stage5_c110_c_ha0), .B(stage5_c111_s_ha0), .So(stage6_c111_s_ha0), .Co(stage6_c111_c_ha0));
    HA ha_201(.A(stage5_c111_c_ha0), .B(stage5_c112_s_ha0), .So(stage6_c112_s_ha0), .Co(stage6_c112_c_ha0));
    HA ha_202(.A(stage5_c112_c_ha0), .B(stage4_c112_c_ha0), .So(stage6_c113_s_ha0), .Co(stage6_c113_c_ha0));
    HA ha_203(.A(stage6_c6_c_ha0), .B(stage6_c7_s_ha0), .So(stage7_c7_s_ha0), .Co(stage7_c7_c_ha0));
    HA ha_204(.A(stage6_c7_c_ha0), .B(stage6_c8_s_ha0), .So(stage7_c8_s_ha0), .Co(stage7_c8_c_ha0));
    HA ha_205(.A(stage6_c8_c_ha0), .B(stage6_c9_s_ha0), .So(stage7_c9_s_ha0), .Co(stage7_c9_c_ha0));
    HA ha_206(.A(stage6_c9_c_ha0), .B(stage6_c10_s_ha0), .So(stage7_c10_s_ha0), .Co(stage7_c10_c_ha0));
    HA ha_207(.A(stage6_c10_c_ha0), .B(stage6_c11_s_ha0), .So(stage7_c11_s_ha0), .Co(stage7_c11_c_ha0));
    HA ha_208(.A(stage6_c11_c_ha0), .B(stage6_c12_s_ha0), .So(stage7_c12_s_ha0), .Co(stage7_c12_c_ha0));
    HA ha_209(.A(stage6_c12_c_ha0), .B(stage6_c13_s_ha0), .So(stage7_c13_s_ha0), .Co(stage7_c13_c_ha0));
    HA ha_210(.A(stage6_c13_c_ha0), .B(stage6_c14_s_ha0), .So(stage7_c14_s_ha0), .Co(stage7_c14_c_ha0));
    HA ha_211(.A(stage6_c14_c_ha0), .B(stage6_c15_s_fa0), .So(stage7_c15_s_ha0), .Co(stage7_c15_c_ha0));
    HA ha_212(.A(stage6_c15_c_fa0), .B(stage6_c16_s_fa0), .So(stage7_c16_s_ha0), .Co(stage7_c16_c_ha0));
    HA ha_213(.A(stage6_c16_c_fa0), .B(stage6_c17_s_fa0), .So(stage7_c17_s_ha0), .Co(stage7_c17_c_ha0));
    HA ha_214(.A(stage6_c17_c_fa0), .B(stage6_c18_s_fa0), .So(stage7_c18_s_ha0), .Co(stage7_c18_c_ha0));
    HA ha_215(.A(stage6_c18_c_fa0), .B(stage6_c19_s_fa0), .So(stage7_c19_s_ha0), .Co(stage7_c19_c_ha0));
    HA ha_216(.A(stage6_c19_c_fa0), .B(stage6_c20_s_fa0), .So(stage7_c20_s_ha0), .Co(stage7_c20_c_ha0));
    HA ha_217(.A(stage6_c20_c_fa0), .B(stage6_c21_s_fa0), .So(stage7_c21_s_ha0), .Co(stage7_c21_c_ha0));
    FA fa_2602(.A(stage6_c21_c_fa0), .B(stage6_c22_s_fa0), .C(stage5_c22_s_ha0), .So(stage7_c22_s_fa0), .Co(stage7_c22_c_fa0));
    FA fa_2603(.A(stage6_c22_c_fa0), .B(stage6_c23_s_fa0), .C(stage5_c23_s_ha0), .So(stage7_c23_s_fa0), .Co(stage7_c23_c_fa0));
    FA fa_2604(.A(stage6_c23_c_fa0), .B(stage6_c24_s_fa0), .C(stage5_c24_s_ha0), .So(stage7_c24_s_fa0), .Co(stage7_c24_c_fa0));
    FA fa_2605(.A(stage6_c24_c_fa0), .B(stage6_c25_s_fa0), .C(stage5_c25_s_fa1), .So(stage7_c25_s_fa0), .Co(stage7_c25_c_fa0));
    FA fa_2606(.A(stage6_c25_c_fa0), .B(stage6_c26_s_fa0), .C(stage5_c26_s_fa1), .So(stage7_c26_s_fa0), .Co(stage7_c26_c_fa0));
    FA fa_2607(.A(stage6_c26_c_fa0), .B(stage6_c27_s_fa0), .C(stage5_c27_s_fa1), .So(stage7_c27_s_fa0), .Co(stage7_c27_c_fa0));
    FA fa_2608(.A(stage6_c27_c_fa0), .B(stage6_c28_s_fa0), .C(stage5_c28_s_fa1), .So(stage7_c28_s_fa0), .Co(stage7_c28_c_fa0));
    FA fa_2609(.A(stage6_c28_c_fa0), .B(stage6_c29_s_fa0), .C(stage5_c29_s_fa1), .So(stage7_c29_s_fa0), .Co(stage7_c29_c_fa0));
    FA fa_2610(.A(stage6_c29_c_fa0), .B(stage6_c30_s_fa0), .C(stage5_c30_s_fa1), .So(stage7_c30_s_fa0), .Co(stage7_c30_c_fa0));
    FA fa_2611(.A(stage6_c30_c_fa0), .B(stage6_c31_s_fa0), .C(stage6_c31_s_ha0), .So(stage7_c31_s_fa0), .Co(stage7_c31_c_fa0));
    FA fa_2612(.A(stage6_c31_c_fa0), .B(stage6_c31_c_ha0), .C(stage6_c32_s_fa0), .So(stage7_c32_s_fa0), .Co(stage7_c32_c_fa0));
    FA fa_2613(.A(stage6_c32_c_fa0), .B(stage6_c32_c_ha0), .C(stage6_c33_s_fa0), .So(stage7_c33_s_fa0), .Co(stage7_c33_c_fa0));
    FA fa_2614(.A(stage6_c33_c_fa0), .B(stage6_c33_c_ha0), .C(stage6_c34_s_fa0), .So(stage7_c34_s_fa0), .Co(stage7_c34_c_fa0));
    FA fa_2615(.A(stage6_c34_c_fa0), .B(stage6_c34_c_ha0), .C(stage6_c35_s_fa0), .So(stage7_c35_s_fa0), .Co(stage7_c35_c_fa0));
    FA fa_2616(.A(stage6_c35_c_fa0), .B(stage6_c35_c_ha0), .C(stage6_c36_s_fa0), .So(stage7_c36_s_fa0), .Co(stage7_c36_c_fa0));
    FA fa_2617(.A(stage6_c36_c_fa0), .B(stage6_c36_c_fa1), .C(stage6_c37_s_fa0), .So(stage7_c37_s_fa0), .Co(stage7_c37_c_fa0));
    FA fa_2618(.A(stage6_c37_c_fa0), .B(stage6_c37_c_fa1), .C(stage6_c38_s_fa0), .So(stage7_c38_s_fa0), .Co(stage7_c38_c_fa0));
    FA fa_2619(.A(stage6_c38_c_fa0), .B(stage6_c38_c_fa1), .C(stage6_c39_s_fa0), .So(stage7_c39_s_fa0), .Co(stage7_c39_c_fa0));
    FA fa_2620(.A(stage6_c39_c_fa0), .B(stage6_c39_c_fa1), .C(stage6_c40_s_fa0), .So(stage7_c40_s_fa0), .Co(stage7_c40_c_fa0));
    FA fa_2621(.A(stage6_c40_c_fa0), .B(stage6_c40_c_fa1), .C(stage6_c41_s_fa0), .So(stage7_c41_s_fa0), .Co(stage7_c41_c_fa0));
    FA fa_2622(.A(stage6_c41_c_fa0), .B(stage6_c41_c_fa1), .C(stage6_c42_s_fa0), .So(stage7_c42_s_fa0), .Co(stage7_c42_c_fa0));
    FA fa_2623(.A(stage6_c42_c_fa0), .B(stage6_c42_c_fa1), .C(stage6_c43_s_fa0), .So(stage7_c43_s_fa0), .Co(stage7_c43_c_fa0));
    FA fa_2624(.A(stage6_c43_c_fa0), .B(stage6_c43_c_fa1), .C(stage6_c44_s_fa0), .So(stage7_c44_s_fa0), .Co(stage7_c44_c_fa0));
    FA fa_2625(.A(stage6_c44_c_fa0), .B(stage6_c44_c_fa1), .C(stage6_c45_s_fa0), .So(stage7_c45_s_fa0), .Co(stage7_c45_c_fa0));
    FA fa_2626(.A(stage6_c45_c_fa0), .B(stage6_c45_c_fa1), .C(stage6_c46_s_fa0), .So(stage7_c46_s_fa0), .Co(stage7_c46_c_fa0));
    FA fa_2627(.A(stage6_c46_c_fa0), .B(stage6_c46_c_fa1), .C(stage6_c47_s_fa0), .So(stage7_c47_s_fa0), .Co(stage7_c47_c_fa0));
    FA fa_2628(.A(stage6_c47_c_fa0), .B(stage6_c47_c_fa1), .C(stage6_c48_s_fa0), .So(stage7_c48_s_fa0), .Co(stage7_c48_c_fa0));
    FA fa_2629(.A(stage6_c48_c_fa0), .B(stage6_c48_c_fa1), .C(stage6_c49_s_fa0), .So(stage7_c49_s_fa0), .Co(stage7_c49_c_fa0));
    FA fa_2630(.A(stage6_c49_c_fa0), .B(stage6_c49_c_fa1), .C(stage6_c50_s_fa0), .So(stage7_c50_s_fa0), .Co(stage7_c50_c_fa0));
    FA fa_2631(.A(stage6_c50_c_fa0), .B(stage6_c50_c_fa1), .C(stage6_c51_s_fa0), .So(stage7_c51_s_fa0), .Co(stage7_c51_c_fa0));
    FA fa_2632(.A(stage6_c51_c_fa0), .B(stage6_c51_c_fa1), .C(stage6_c52_s_fa0), .So(stage7_c52_s_fa0), .Co(stage7_c52_c_fa0));
    FA fa_2633(.A(stage6_c52_c_fa0), .B(stage6_c52_c_fa1), .C(stage6_c53_s_fa0), .So(stage7_c53_s_fa0), .Co(stage7_c53_c_fa0));
    FA fa_2634(.A(stage6_c53_c_fa0), .B(stage6_c53_c_fa1), .C(stage6_c54_s_fa0), .So(stage7_c54_s_fa0), .Co(stage7_c54_c_fa0));
    FA fa_2635(.A(stage6_c54_c_fa0), .B(stage6_c54_c_fa1), .C(stage6_c55_s_fa0), .So(stage7_c55_s_fa0), .Co(stage7_c55_c_fa0));
    FA fa_2636(.A(stage6_c55_c_fa0), .B(stage6_c55_c_fa1), .C(stage6_c56_s_fa0), .So(stage7_c56_s_fa0), .Co(stage7_c56_c_fa0));
    FA fa_2637(.A(stage6_c56_c_fa0), .B(stage6_c56_c_fa1), .C(stage6_c57_s_fa0), .So(stage7_c57_s_fa0), .Co(stage7_c57_c_fa0));
    FA fa_2638(.A(stage6_c57_c_fa0), .B(stage6_c57_c_fa1), .C(stage6_c58_s_fa0), .So(stage7_c58_s_fa0), .Co(stage7_c58_c_fa0));
    FA fa_2639(.A(stage6_c58_c_fa0), .B(stage6_c58_c_fa1), .C(stage6_c59_s_fa0), .So(stage7_c59_s_fa0), .Co(stage7_c59_c_fa0));
    FA fa_2640(.A(stage6_c59_c_fa0), .B(stage6_c59_c_fa1), .C(stage6_c60_s_fa0), .So(stage7_c60_s_fa0), .Co(stage7_c60_c_fa0));
    FA fa_2641(.A(stage6_c60_c_fa0), .B(stage6_c60_c_fa1), .C(stage6_c61_s_fa0), .So(stage7_c61_s_fa0), .Co(stage7_c61_c_fa0));
    FA fa_2642(.A(stage6_c61_c_fa0), .B(stage6_c61_c_fa1), .C(stage6_c62_s_fa0), .So(stage7_c62_s_fa0), .Co(stage7_c62_c_fa0));
    FA fa_2643(.A(stage6_c62_c_fa0), .B(stage6_c62_c_fa1), .C(stage6_c63_s_fa0), .So(stage7_c63_s_fa0), .Co(stage7_c63_c_fa0));
    FA fa_2644(.A(stage6_c63_c_fa0), .B(stage6_c63_c_fa1), .C(stage6_c64_s_fa0), .So(stage7_c64_s_fa0), .Co(stage7_c64_c_fa0));
    FA fa_2645(.A(stage6_c64_c_fa0), .B(stage6_c64_c_fa1), .C(stage6_c65_s_fa0), .So(stage7_c65_s_fa0), .Co(stage7_c65_c_fa0));
    FA fa_2646(.A(stage6_c65_c_fa0), .B(stage6_c65_c_fa1), .C(stage6_c66_s_fa0), .So(stage7_c66_s_fa0), .Co(stage7_c66_c_fa0));
    FA fa_2647(.A(stage6_c66_c_fa0), .B(stage6_c66_c_fa1), .C(stage6_c67_s_fa0), .So(stage7_c67_s_fa0), .Co(stage7_c67_c_fa0));
    FA fa_2648(.A(stage6_c67_c_fa0), .B(stage6_c67_c_fa1), .C(stage6_c68_s_fa0), .So(stage7_c68_s_fa0), .Co(stage7_c68_c_fa0));
    FA fa_2649(.A(stage6_c68_c_fa0), .B(stage6_c68_c_fa1), .C(stage6_c69_s_fa0), .So(stage7_c69_s_fa0), .Co(stage7_c69_c_fa0));
    FA fa_2650(.A(stage6_c69_c_fa0), .B(stage6_c69_c_fa1), .C(stage6_c70_s_fa0), .So(stage7_c70_s_fa0), .Co(stage7_c70_c_fa0));
    FA fa_2651(.A(stage6_c70_c_fa0), .B(stage6_c70_c_fa1), .C(stage6_c71_s_fa0), .So(stage7_c71_s_fa0), .Co(stage7_c71_c_fa0));
    FA fa_2652(.A(stage6_c71_c_fa0), .B(stage6_c71_c_fa1), .C(stage6_c72_s_fa0), .So(stage7_c72_s_fa0), .Co(stage7_c72_c_fa0));
    FA fa_2653(.A(stage6_c72_c_fa0), .B(stage6_c72_c_fa1), .C(stage6_c73_s_fa0), .So(stage7_c73_s_fa0), .Co(stage7_c73_c_fa0));
    FA fa_2654(.A(stage6_c73_c_fa0), .B(stage6_c73_c_fa1), .C(stage6_c74_s_fa0), .So(stage7_c74_s_fa0), .Co(stage7_c74_c_fa0));
    FA fa_2655(.A(stage6_c74_c_fa0), .B(stage6_c74_c_fa1), .C(stage6_c75_s_fa0), .So(stage7_c75_s_fa0), .Co(stage7_c75_c_fa0));
    FA fa_2656(.A(stage6_c75_c_fa0), .B(stage6_c75_c_fa1), .C(stage6_c76_s_fa0), .So(stage7_c76_s_fa0), .Co(stage7_c76_c_fa0));
    FA fa_2657(.A(stage6_c76_c_fa0), .B(stage6_c76_c_fa1), .C(stage6_c77_s_fa0), .So(stage7_c77_s_fa0), .Co(stage7_c77_c_fa0));
    FA fa_2658(.A(stage6_c77_c_fa0), .B(stage6_c77_c_fa1), .C(stage6_c78_s_fa0), .So(stage7_c78_s_fa0), .Co(stage7_c78_c_fa0));
    FA fa_2659(.A(stage6_c78_c_fa0), .B(stage6_c78_c_fa1), .C(stage6_c79_s_fa0), .So(stage7_c79_s_fa0), .Co(stage7_c79_c_fa0));
    FA fa_2660(.A(stage6_c79_c_fa0), .B(stage6_c79_c_fa1), .C(stage6_c80_s_fa0), .So(stage7_c80_s_fa0), .Co(stage7_c80_c_fa0));
    FA fa_2661(.A(stage6_c80_c_fa0), .B(stage6_c80_c_fa1), .C(stage6_c81_s_fa0), .So(stage7_c81_s_fa0), .Co(stage7_c81_c_fa0));
    FA fa_2662(.A(stage6_c81_c_fa0), .B(stage6_c81_c_fa1), .C(stage6_c82_s_fa0), .So(stage7_c82_s_fa0), .Co(stage7_c82_c_fa0));
    FA fa_2663(.A(stage6_c82_c_fa0), .B(stage6_c82_c_ha0), .C(stage6_c83_s_fa0), .So(stage7_c83_s_fa0), .Co(stage7_c83_c_fa0));
    FA fa_2664(.A(stage6_c83_c_fa0), .B(stage6_c83_c_ha0), .C(stage6_c84_s_fa0), .So(stage7_c84_s_fa0), .Co(stage7_c84_c_fa0));
    FA fa_2665(.A(stage6_c84_c_fa0), .B(stage6_c84_c_ha0), .C(stage6_c85_s_fa0), .So(stage7_c85_s_fa0), .Co(stage7_c85_c_fa0));
    FA fa_2666(.A(stage6_c85_c_fa0), .B(stage6_c85_c_ha0), .C(stage6_c86_s_fa0), .So(stage7_c86_s_fa0), .Co(stage7_c86_c_fa0));
    FA fa_2667(.A(stage6_c86_c_fa0), .B(stage6_c87_s_fa0), .C(stage5_c87_s_fa1), .So(stage7_c87_s_fa0), .Co(stage7_c87_c_fa0));
    FA fa_2668(.A(stage6_c87_c_fa0), .B(stage6_c88_s_fa0), .C(stage5_c88_s_fa1), .So(stage7_c88_s_fa0), .Co(stage7_c88_c_fa0));
    FA fa_2669(.A(stage6_c88_c_fa0), .B(stage6_c89_s_fa0), .C(stage5_c89_s_fa1), .So(stage7_c89_s_fa0), .Co(stage7_c89_c_fa0));
    FA fa_2670(.A(stage6_c89_c_fa0), .B(stage6_c90_s_fa0), .C(stage5_c90_s_fa1), .So(stage7_c90_s_fa0), .Co(stage7_c90_c_fa0));
    FA fa_2671(.A(stage6_c90_c_fa0), .B(stage6_c91_s_fa0), .C(stage5_c91_s_fa1), .So(stage7_c91_s_fa0), .Co(stage7_c91_c_fa0));
    FA fa_2672(.A(stage6_c91_c_fa0), .B(stage6_c92_s_fa0), .C(stage5_c92_s_fa1), .So(stage7_c92_s_fa0), .Co(stage7_c92_c_fa0));
    FA fa_2673(.A(stage6_c92_c_fa0), .B(stage6_c93_s_fa0), .C(stage5_c93_s_ha0), .So(stage7_c93_s_fa0), .Co(stage7_c93_c_fa0));
    FA fa_2674(.A(stage6_c93_c_fa0), .B(stage6_c94_s_fa0), .C(stage4_c94_s_fa1), .So(stage7_c94_s_fa0), .Co(stage7_c94_c_fa0));
    HA ha_218(.A(stage6_c94_c_fa0), .B(stage6_c95_s_fa0), .So(stage7_c95_s_ha0), .Co(stage7_c95_c_ha0));
    HA ha_219(.A(stage6_c95_c_fa0), .B(stage6_c96_s_fa0), .So(stage7_c96_s_ha0), .Co(stage7_c96_c_ha0));
    HA ha_220(.A(stage6_c96_c_fa0), .B(stage6_c97_s_fa0), .So(stage7_c97_s_ha0), .Co(stage7_c97_c_ha0));
    HA ha_221(.A(stage6_c97_c_fa0), .B(stage6_c98_s_fa0), .So(stage7_c98_s_ha0), .Co(stage7_c98_c_ha0));
    HA ha_222(.A(stage6_c98_c_fa0), .B(stage6_c99_s_fa0), .So(stage7_c99_s_ha0), .Co(stage7_c99_c_ha0));
    HA ha_223(.A(stage6_c99_c_fa0), .B(stage6_c100_s_fa0), .So(stage7_c100_s_ha0), .Co(stage7_c100_c_ha0));
    HA ha_224(.A(stage6_c100_c_fa0), .B(stage6_c101_s_ha0), .So(stage7_c101_s_ha0), .Co(stage7_c101_c_ha0));
    HA ha_225(.A(stage6_c101_c_ha0), .B(stage6_c102_s_ha0), .So(stage7_c102_s_ha0), .Co(stage7_c102_c_ha0));
    HA ha_226(.A(stage6_c102_c_ha0), .B(stage6_c103_s_ha0), .So(stage7_c103_s_ha0), .Co(stage7_c103_c_ha0));
    HA ha_227(.A(stage6_c103_c_ha0), .B(stage6_c104_s_ha0), .So(stage7_c104_s_ha0), .Co(stage7_c104_c_ha0));
    HA ha_228(.A(stage6_c104_c_ha0), .B(stage6_c105_s_ha0), .So(stage7_c105_s_ha0), .Co(stage7_c105_c_ha0));
    HA ha_229(.A(stage6_c105_c_ha0), .B(stage6_c106_s_ha0), .So(stage7_c106_s_ha0), .Co(stage7_c106_c_ha0));
    HA ha_230(.A(stage6_c106_c_ha0), .B(stage6_c107_s_ha0), .So(stage7_c107_s_ha0), .Co(stage7_c107_c_ha0));
    HA ha_231(.A(stage6_c107_c_ha0), .B(stage6_c108_s_ha0), .So(stage7_c108_s_ha0), .Co(stage7_c108_c_ha0));
    HA ha_232(.A(stage6_c108_c_ha0), .B(stage6_c109_s_ha0), .So(stage7_c109_s_ha0), .Co(stage7_c109_c_ha0));
    HA ha_233(.A(stage6_c109_c_ha0), .B(stage6_c110_s_ha0), .So(stage7_c110_s_ha0), .Co(stage7_c110_c_ha0));
    HA ha_234(.A(stage6_c110_c_ha0), .B(stage6_c111_s_ha0), .So(stage7_c111_s_ha0), .Co(stage7_c111_c_ha0));
    HA ha_235(.A(stage6_c111_c_ha0), .B(stage6_c112_s_ha0), .So(stage7_c112_s_ha0), .Co(stage7_c112_c_ha0));
    HA ha_236(.A(stage6_c112_c_ha0), .B(stage6_c113_s_ha0), .So(stage7_c113_s_ha0), .Co(stage7_c113_c_ha0));
    HA ha_237(.A(stage7_c7_c_ha0), .B(stage7_c8_s_ha0), .So(stage8_c8_s_ha0), .Co(stage8_c8_c_ha0));
    HA ha_238(.A(stage7_c8_c_ha0), .B(stage7_c9_s_ha0), .So(stage8_c9_s_ha0), .Co(stage8_c9_c_ha0));
    HA ha_239(.A(stage7_c9_c_ha0), .B(stage7_c10_s_ha0), .So(stage8_c10_s_ha0), .Co(stage8_c10_c_ha0));
    HA ha_240(.A(stage7_c10_c_ha0), .B(stage7_c11_s_ha0), .So(stage8_c11_s_ha0), .Co(stage8_c11_c_ha0));
    HA ha_241(.A(stage7_c11_c_ha0), .B(stage7_c12_s_ha0), .So(stage8_c12_s_ha0), .Co(stage8_c12_c_ha0));
    HA ha_242(.A(stage7_c12_c_ha0), .B(stage7_c13_s_ha0), .So(stage8_c13_s_ha0), .Co(stage8_c13_c_ha0));
    HA ha_243(.A(stage7_c13_c_ha0), .B(stage7_c14_s_ha0), .So(stage8_c14_s_ha0), .Co(stage8_c14_c_ha0));
    HA ha_244(.A(stage7_c14_c_ha0), .B(stage7_c15_s_ha0), .So(stage8_c15_s_ha0), .Co(stage8_c15_c_ha0));
    HA ha_245(.A(stage7_c15_c_ha0), .B(stage7_c16_s_ha0), .So(stage8_c16_s_ha0), .Co(stage8_c16_c_ha0));
    HA ha_246(.A(stage7_c16_c_ha0), .B(stage7_c17_s_ha0), .So(stage8_c17_s_ha0), .Co(stage8_c17_c_ha0));
    HA ha_247(.A(stage7_c17_c_ha0), .B(stage7_c18_s_ha0), .So(stage8_c18_s_ha0), .Co(stage8_c18_c_ha0));
    HA ha_248(.A(stage7_c18_c_ha0), .B(stage7_c19_s_ha0), .So(stage8_c19_s_ha0), .Co(stage8_c19_c_ha0));
    HA ha_249(.A(stage7_c19_c_ha0), .B(stage7_c20_s_ha0), .So(stage8_c20_s_ha0), .Co(stage8_c20_c_ha0));
    HA ha_250(.A(stage7_c20_c_ha0), .B(stage7_c21_s_ha0), .So(stage8_c21_s_ha0), .Co(stage8_c21_c_ha0));
    HA ha_251(.A(stage7_c21_c_ha0), .B(stage7_c22_s_fa0), .So(stage8_c22_s_ha0), .Co(stage8_c22_c_ha0));
    HA ha_252(.A(stage7_c22_c_fa0), .B(stage7_c23_s_fa0), .So(stage8_c23_s_ha0), .Co(stage8_c23_c_ha0));
    HA ha_253(.A(stage7_c23_c_fa0), .B(stage7_c24_s_fa0), .So(stage8_c24_s_ha0), .Co(stage8_c24_c_ha0));
    HA ha_254(.A(stage7_c24_c_fa0), .B(stage7_c25_s_fa0), .So(stage8_c25_s_ha0), .Co(stage8_c25_c_ha0));
    HA ha_255(.A(stage7_c25_c_fa0), .B(stage7_c26_s_fa0), .So(stage8_c26_s_ha0), .Co(stage8_c26_c_ha0));
    HA ha_256(.A(stage7_c26_c_fa0), .B(stage7_c27_s_fa0), .So(stage8_c27_s_ha0), .Co(stage8_c27_c_ha0));
    HA ha_257(.A(stage7_c27_c_fa0), .B(stage7_c28_s_fa0), .So(stage8_c28_s_ha0), .Co(stage8_c28_c_ha0));
    HA ha_258(.A(stage7_c28_c_fa0), .B(stage7_c29_s_fa0), .So(stage8_c29_s_ha0), .Co(stage8_c29_c_ha0));
    HA ha_259(.A(stage7_c29_c_fa0), .B(stage7_c30_s_fa0), .So(stage8_c30_s_ha0), .Co(stage8_c30_c_ha0));
    HA ha_260(.A(stage7_c30_c_fa0), .B(stage7_c31_s_fa0), .So(stage8_c31_s_ha0), .Co(stage8_c31_c_ha0));
    FA fa_2675(.A(stage7_c31_c_fa0), .B(stage7_c32_s_fa0), .C(stage6_c32_s_ha0), .So(stage8_c32_s_fa0), .Co(stage8_c32_c_fa0));
    FA fa_2676(.A(stage7_c32_c_fa0), .B(stage7_c33_s_fa0), .C(stage6_c33_s_ha0), .So(stage8_c33_s_fa0), .Co(stage8_c33_c_fa0));
    FA fa_2677(.A(stage7_c33_c_fa0), .B(stage7_c34_s_fa0), .C(stage6_c34_s_ha0), .So(stage8_c34_s_fa0), .Co(stage8_c34_c_fa0));
    FA fa_2678(.A(stage7_c34_c_fa0), .B(stage7_c35_s_fa0), .C(stage6_c35_s_ha0), .So(stage8_c35_s_fa0), .Co(stage8_c35_c_fa0));
    FA fa_2679(.A(stage7_c35_c_fa0), .B(stage7_c36_s_fa0), .C(stage6_c36_s_fa1), .So(stage8_c36_s_fa0), .Co(stage8_c36_c_fa0));
    FA fa_2680(.A(stage7_c36_c_fa0), .B(stage7_c37_s_fa0), .C(stage6_c37_s_fa1), .So(stage8_c37_s_fa0), .Co(stage8_c37_c_fa0));
    FA fa_2681(.A(stage7_c37_c_fa0), .B(stage7_c38_s_fa0), .C(stage6_c38_s_fa1), .So(stage8_c38_s_fa0), .Co(stage8_c38_c_fa0));
    FA fa_2682(.A(stage7_c38_c_fa0), .B(stage7_c39_s_fa0), .C(stage6_c39_s_fa1), .So(stage8_c39_s_fa0), .Co(stage8_c39_c_fa0));
    FA fa_2683(.A(stage7_c39_c_fa0), .B(stage7_c40_s_fa0), .C(stage6_c40_s_fa1), .So(stage8_c40_s_fa0), .Co(stage8_c40_c_fa0));
    FA fa_2684(.A(stage7_c40_c_fa0), .B(stage7_c41_s_fa0), .C(stage6_c41_s_fa1), .So(stage8_c41_s_fa0), .Co(stage8_c41_c_fa0));
    FA fa_2685(.A(stage7_c41_c_fa0), .B(stage7_c42_s_fa0), .C(stage6_c42_s_fa1), .So(stage8_c42_s_fa0), .Co(stage8_c42_c_fa0));
    FA fa_2686(.A(stage7_c42_c_fa0), .B(stage7_c43_s_fa0), .C(stage6_c43_s_fa1), .So(stage8_c43_s_fa0), .Co(stage8_c43_c_fa0));
    FA fa_2687(.A(stage7_c43_c_fa0), .B(stage7_c44_s_fa0), .C(stage6_c44_s_fa1), .So(stage8_c44_s_fa0), .Co(stage8_c44_c_fa0));
    FA fa_2688(.A(stage7_c44_c_fa0), .B(stage7_c45_s_fa0), .C(stage6_c45_s_fa1), .So(stage8_c45_s_fa0), .Co(stage8_c45_c_fa0));
    FA fa_2689(.A(stage7_c45_c_fa0), .B(stage7_c46_s_fa0), .C(stage6_c46_s_fa1), .So(stage8_c46_s_fa0), .Co(stage8_c46_c_fa0));
    FA fa_2690(.A(stage7_c46_c_fa0), .B(stage7_c47_s_fa0), .C(stage6_c47_s_fa1), .So(stage8_c47_s_fa0), .Co(stage8_c47_c_fa0));
    FA fa_2691(.A(stage7_c47_c_fa0), .B(stage7_c48_s_fa0), .C(stage6_c48_s_fa1), .So(stage8_c48_s_fa0), .Co(stage8_c48_c_fa0));
    FA fa_2692(.A(stage7_c48_c_fa0), .B(stage7_c49_s_fa0), .C(stage6_c49_s_fa1), .So(stage8_c49_s_fa0), .Co(stage8_c49_c_fa0));
    FA fa_2693(.A(stage7_c49_c_fa0), .B(stage7_c50_s_fa0), .C(stage6_c50_s_fa1), .So(stage8_c50_s_fa0), .Co(stage8_c50_c_fa0));
    FA fa_2694(.A(stage7_c50_c_fa0), .B(stage7_c51_s_fa0), .C(stage6_c51_s_fa1), .So(stage8_c51_s_fa0), .Co(stage8_c51_c_fa0));
    FA fa_2695(.A(stage7_c51_c_fa0), .B(stage7_c52_s_fa0), .C(stage6_c52_s_fa1), .So(stage8_c52_s_fa0), .Co(stage8_c52_c_fa0));
    FA fa_2696(.A(stage7_c52_c_fa0), .B(stage7_c53_s_fa0), .C(stage6_c53_s_fa1), .So(stage8_c53_s_fa0), .Co(stage8_c53_c_fa0));
    FA fa_2697(.A(stage7_c53_c_fa0), .B(stage7_c54_s_fa0), .C(stage6_c54_s_fa1), .So(stage8_c54_s_fa0), .Co(stage8_c54_c_fa0));
    FA fa_2698(.A(stage7_c54_c_fa0), .B(stage7_c55_s_fa0), .C(stage6_c55_s_fa1), .So(stage8_c55_s_fa0), .Co(stage8_c55_c_fa0));
    FA fa_2699(.A(stage7_c55_c_fa0), .B(stage7_c56_s_fa0), .C(stage6_c56_s_fa1), .So(stage8_c56_s_fa0), .Co(stage8_c56_c_fa0));
    FA fa_2700(.A(stage7_c56_c_fa0), .B(stage7_c57_s_fa0), .C(stage6_c57_s_fa1), .So(stage8_c57_s_fa0), .Co(stage8_c57_c_fa0));
    FA fa_2701(.A(stage7_c57_c_fa0), .B(stage7_c58_s_fa0), .C(stage6_c58_s_fa1), .So(stage8_c58_s_fa0), .Co(stage8_c58_c_fa0));
    FA fa_2702(.A(stage7_c58_c_fa0), .B(stage7_c59_s_fa0), .C(stage6_c59_s_fa1), .So(stage8_c59_s_fa0), .Co(stage8_c59_c_fa0));
    FA fa_2703(.A(stage7_c59_c_fa0), .B(stage7_c60_s_fa0), .C(stage6_c60_s_fa1), .So(stage8_c60_s_fa0), .Co(stage8_c60_c_fa0));
    FA fa_2704(.A(stage7_c60_c_fa0), .B(stage7_c61_s_fa0), .C(stage6_c61_s_fa1), .So(stage8_c61_s_fa0), .Co(stage8_c61_c_fa0));
    FA fa_2705(.A(stage7_c61_c_fa0), .B(stage7_c62_s_fa0), .C(stage6_c62_s_fa1), .So(stage8_c62_s_fa0), .Co(stage8_c62_c_fa0));
    FA fa_2706(.A(stage7_c62_c_fa0), .B(stage7_c63_s_fa0), .C(stage6_c63_s_fa1), .So(stage8_c63_s_fa0), .Co(stage8_c63_c_fa0));
    FA fa_2707(.A(stage7_c63_c_fa0), .B(stage7_c64_s_fa0), .C(stage6_c64_s_fa1), .So(stage8_c64_s_fa0), .Co(stage8_c64_c_fa0));
    FA fa_2708(.A(stage7_c64_c_fa0), .B(stage7_c65_s_fa0), .C(stage6_c65_s_fa1), .So(stage8_c65_s_fa0), .Co(stage8_c65_c_fa0));
    FA fa_2709(.A(stage7_c65_c_fa0), .B(stage7_c66_s_fa0), .C(stage6_c66_s_fa1), .So(stage8_c66_s_fa0), .Co(stage8_c66_c_fa0));
    FA fa_2710(.A(stage7_c66_c_fa0), .B(stage7_c67_s_fa0), .C(stage6_c67_s_fa1), .So(stage8_c67_s_fa0), .Co(stage8_c67_c_fa0));
    FA fa_2711(.A(stage7_c67_c_fa0), .B(stage7_c68_s_fa0), .C(stage6_c68_s_fa1), .So(stage8_c68_s_fa0), .Co(stage8_c68_c_fa0));
    FA fa_2712(.A(stage7_c68_c_fa0), .B(stage7_c69_s_fa0), .C(stage6_c69_s_fa1), .So(stage8_c69_s_fa0), .Co(stage8_c69_c_fa0));
    FA fa_2713(.A(stage7_c69_c_fa0), .B(stage7_c70_s_fa0), .C(stage6_c70_s_fa1), .So(stage8_c70_s_fa0), .Co(stage8_c70_c_fa0));
    FA fa_2714(.A(stage7_c70_c_fa0), .B(stage7_c71_s_fa0), .C(stage6_c71_s_fa1), .So(stage8_c71_s_fa0), .Co(stage8_c71_c_fa0));
    FA fa_2715(.A(stage7_c71_c_fa0), .B(stage7_c72_s_fa0), .C(stage6_c72_s_fa1), .So(stage8_c72_s_fa0), .Co(stage8_c72_c_fa0));
    FA fa_2716(.A(stage7_c72_c_fa0), .B(stage7_c73_s_fa0), .C(stage6_c73_s_fa1), .So(stage8_c73_s_fa0), .Co(stage8_c73_c_fa0));
    FA fa_2717(.A(stage7_c73_c_fa0), .B(stage7_c74_s_fa0), .C(stage6_c74_s_fa1), .So(stage8_c74_s_fa0), .Co(stage8_c74_c_fa0));
    FA fa_2718(.A(stage7_c74_c_fa0), .B(stage7_c75_s_fa0), .C(stage6_c75_s_fa1), .So(stage8_c75_s_fa0), .Co(stage8_c75_c_fa0));
    FA fa_2719(.A(stage7_c75_c_fa0), .B(stage7_c76_s_fa0), .C(stage6_c76_s_fa1), .So(stage8_c76_s_fa0), .Co(stage8_c76_c_fa0));
    FA fa_2720(.A(stage7_c76_c_fa0), .B(stage7_c77_s_fa0), .C(stage6_c77_s_fa1), .So(stage8_c77_s_fa0), .Co(stage8_c77_c_fa0));
    FA fa_2721(.A(stage7_c77_c_fa0), .B(stage7_c78_s_fa0), .C(stage6_c78_s_fa1), .So(stage8_c78_s_fa0), .Co(stage8_c78_c_fa0));
    FA fa_2722(.A(stage7_c78_c_fa0), .B(stage7_c79_s_fa0), .C(stage6_c79_s_fa1), .So(stage8_c79_s_fa0), .Co(stage8_c79_c_fa0));
    FA fa_2723(.A(stage7_c79_c_fa0), .B(stage7_c80_s_fa0), .C(stage6_c80_s_fa1), .So(stage8_c80_s_fa0), .Co(stage8_c80_c_fa0));
    FA fa_2724(.A(stage7_c80_c_fa0), .B(stage7_c81_s_fa0), .C(stage6_c81_s_fa1), .So(stage8_c81_s_fa0), .Co(stage8_c81_c_fa0));
    FA fa_2725(.A(stage7_c81_c_fa0), .B(stage7_c82_s_fa0), .C(stage6_c82_s_ha0), .So(stage8_c82_s_fa0), .Co(stage8_c82_c_fa0));
    FA fa_2726(.A(stage7_c82_c_fa0), .B(stage7_c83_s_fa0), .C(stage6_c83_s_ha0), .So(stage8_c83_s_fa0), .Co(stage8_c83_c_fa0));
    FA fa_2727(.A(stage7_c83_c_fa0), .B(stage7_c84_s_fa0), .C(stage6_c84_s_ha0), .So(stage8_c84_s_fa0), .Co(stage8_c84_c_fa0));
    FA fa_2728(.A(stage7_c84_c_fa0), .B(stage7_c85_s_fa0), .C(stage6_c85_s_ha0), .So(stage8_c85_s_fa0), .Co(stage8_c85_c_fa0));
    FA fa_2729(.A(stage7_c85_c_fa0), .B(stage7_c86_s_fa0), .C(stage5_c86_s_fa1), .So(stage8_c86_s_fa0), .Co(stage8_c86_c_fa0));
    HA ha_261(.A(stage7_c86_c_fa0), .B(stage7_c87_s_fa0), .So(stage8_c87_s_ha0), .Co(stage8_c87_c_ha0));
    HA ha_262(.A(stage7_c87_c_fa0), .B(stage7_c88_s_fa0), .So(stage8_c88_s_ha0), .Co(stage8_c88_c_ha0));
    HA ha_263(.A(stage7_c88_c_fa0), .B(stage7_c89_s_fa0), .So(stage8_c89_s_ha0), .Co(stage8_c89_c_ha0));
    HA ha_264(.A(stage7_c89_c_fa0), .B(stage7_c90_s_fa0), .So(stage8_c90_s_ha0), .Co(stage8_c90_c_ha0));
    HA ha_265(.A(stage7_c90_c_fa0), .B(stage7_c91_s_fa0), .So(stage8_c91_s_ha0), .Co(stage8_c91_c_ha0));
    HA ha_266(.A(stage7_c91_c_fa0), .B(stage7_c92_s_fa0), .So(stage8_c92_s_ha0), .Co(stage8_c92_c_ha0));
    HA ha_267(.A(stage7_c92_c_fa0), .B(stage7_c93_s_fa0), .So(stage8_c93_s_ha0), .Co(stage8_c93_c_ha0));
    HA ha_268(.A(stage7_c93_c_fa0), .B(stage7_c94_s_fa0), .So(stage8_c94_s_ha0), .Co(stage8_c94_c_ha0));
    HA ha_269(.A(stage7_c94_c_fa0), .B(stage7_c95_s_ha0), .So(stage8_c95_s_ha0), .Co(stage8_c95_c_ha0));
    HA ha_270(.A(stage7_c95_c_ha0), .B(stage7_c96_s_ha0), .So(stage8_c96_s_ha0), .Co(stage8_c96_c_ha0));
    HA ha_271(.A(stage7_c96_c_ha0), .B(stage7_c97_s_ha0), .So(stage8_c97_s_ha0), .Co(stage8_c97_c_ha0));
    HA ha_272(.A(stage7_c97_c_ha0), .B(stage7_c98_s_ha0), .So(stage8_c98_s_ha0), .Co(stage8_c98_c_ha0));
    HA ha_273(.A(stage7_c98_c_ha0), .B(stage7_c99_s_ha0), .So(stage8_c99_s_ha0), .Co(stage8_c99_c_ha0));
    HA ha_274(.A(stage7_c99_c_ha0), .B(stage7_c100_s_ha0), .So(stage8_c100_s_ha0), .Co(stage8_c100_c_ha0));
    HA ha_275(.A(stage7_c100_c_ha0), .B(stage7_c101_s_ha0), .So(stage8_c101_s_ha0), .Co(stage8_c101_c_ha0));
    HA ha_276(.A(stage7_c101_c_ha0), .B(stage7_c102_s_ha0), .So(stage8_c102_s_ha0), .Co(stage8_c102_c_ha0));
    HA ha_277(.A(stage7_c102_c_ha0), .B(stage7_c103_s_ha0), .So(stage8_c103_s_ha0), .Co(stage8_c103_c_ha0));
    HA ha_278(.A(stage7_c103_c_ha0), .B(stage7_c104_s_ha0), .So(stage8_c104_s_ha0), .Co(stage8_c104_c_ha0));
    HA ha_279(.A(stage7_c104_c_ha0), .B(stage7_c105_s_ha0), .So(stage8_c105_s_ha0), .Co(stage8_c105_c_ha0));
    HA ha_280(.A(stage7_c105_c_ha0), .B(stage7_c106_s_ha0), .So(stage8_c106_s_ha0), .Co(stage8_c106_c_ha0));
    HA ha_281(.A(stage7_c106_c_ha0), .B(stage7_c107_s_ha0), .So(stage8_c107_s_ha0), .Co(stage8_c107_c_ha0));
    HA ha_282(.A(stage7_c107_c_ha0), .B(stage7_c108_s_ha0), .So(stage8_c108_s_ha0), .Co(stage8_c108_c_ha0));
    HA ha_283(.A(stage7_c108_c_ha0), .B(stage7_c109_s_ha0), .So(stage8_c109_s_ha0), .Co(stage8_c109_c_ha0));
    HA ha_284(.A(stage7_c109_c_ha0), .B(stage7_c110_s_ha0), .So(stage8_c110_s_ha0), .Co(stage8_c110_c_ha0));
    HA ha_285(.A(stage7_c110_c_ha0), .B(stage7_c111_s_ha0), .So(stage8_c111_s_ha0), .Co(stage8_c111_c_ha0));
    HA ha_286(.A(stage7_c111_c_ha0), .B(stage7_c112_s_ha0), .So(stage8_c112_s_ha0), .Co(stage8_c112_c_ha0));
    HA ha_287(.A(stage7_c112_c_ha0), .B(stage7_c113_s_ha0), .So(stage8_c113_s_ha0), .Co(stage8_c113_c_ha0));
    HA ha_288(.A(stage7_c113_c_ha0), .B(stage6_c113_c_ha0), .So(stage8_c114_s_ha0), .Co(stage8_c114_c_ha0));
endmodule


module HA(A, B, So, Co);
    input A, B;
    output So, Co;

    assign So = A ^ B;
    assign Co = A & B;
endmodule

module FA(A, B, C, So, Co);
    input A, B, C;
    output So, Co;

    assign So = A ^ B ^ C;
    assign Co = (A & B) | (C & (A | B));
endmodule

