



module INVX1 (A, Y);
input  A ;
output Y ;

endmodule



module INVX4 (Y, A);
input  A ;
output Y ;

endmodule



module NAND2X1 (A, B, Y);
input  A ;
input  B ;
output Y ;

endmodule



module NOR2X1 (A, B, Y);
input  A ;
input  B ;
output Y ;

endmodule


